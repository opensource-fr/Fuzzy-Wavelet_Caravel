// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire clknet_0_wb_clk_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _298_ (.I(net242),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _299_ (.I(net206),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _300_ (.A1(net103),
    .A2(net66),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _301_ (.I(_067_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _302_ (.I(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _303_ (.I(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _304_ (.A1(_066_),
    .A2(_070_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _305_ (.A1(_065_),
    .A2(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _306_ (.I(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _307_ (.I(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _308_ (.I(_074_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _309_ (.I(net142),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _310_ (.I(_073_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _311_ (.A1(net207),
    .A2(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _312_ (.A1(_075_),
    .A2(_000_),
    .B(_077_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _313_ (.I0(net218),
    .I1(net153),
    .S(_074_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _314_ (.I(_078_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _315_ (.I0(net229),
    .I1(net164),
    .S(_074_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _316_ (.I(_079_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _317_ (.I0(net232),
    .I1(net167),
    .S(_074_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _318_ (.I(_080_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _319_ (.I0(net233),
    .I1(net168),
    .S(_074_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(_081_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _321_ (.I(_073_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _322_ (.I0(net234),
    .I1(net169),
    .S(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _323_ (.I(_083_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _324_ (.I0(net235),
    .I1(net170),
    .S(_082_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _325_ (.I(_084_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _326_ (.I(net171),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _327_ (.A1(net236),
    .A2(_076_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _328_ (.A1(_085_),
    .A2(_000_),
    .B(_086_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _329_ (.I0(net237),
    .I1(net172),
    .S(_082_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _330_ (.I(_087_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _331_ (.I0(net238),
    .I1(net173),
    .S(_082_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _332_ (.I(_088_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _333_ (.I(net143),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _334_ (.A1(net208),
    .A2(_076_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _335_ (.A1(_089_),
    .A2(_000_),
    .B(_090_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _336_ (.I0(net209),
    .I1(net144),
    .S(_082_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _337_ (.I(_091_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _338_ (.I0(net210),
    .I1(net145),
    .S(_082_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _339_ (.I(_092_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _340_ (.I0(net211),
    .I1(net146),
    .S(_082_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _341_ (.I(_093_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _342_ (.I(net147),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _343_ (.A1(net212),
    .A2(_076_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _344_ (.A1(_094_),
    .A2(_000_),
    .B(_095_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _345_ (.I(net148),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _346_ (.A1(net213),
    .A2(_076_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _347_ (.A1(_096_),
    .A2(_000_),
    .B(_097_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _348_ (.I0(net214),
    .I1(net149),
    .S(_082_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _349_ (.I(_098_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _350_ (.I0(net215),
    .I1(net150),
    .S(_082_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _351_ (.I(_099_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _352_ (.I0(net216),
    .I1(net151),
    .S(_082_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _353_ (.I(_100_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _354_ (.I0(net217),
    .I1(net152),
    .S(_073_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _355_ (.I(_101_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _356_ (.I0(net219),
    .I1(net154),
    .S(_073_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _357_ (.I(_102_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _358_ (.I0(net220),
    .I1(net155),
    .S(_073_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _359_ (.I(_103_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _360_ (.I(net156),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _361_ (.A1(net221),
    .A2(_076_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _362_ (.A1(_104_),
    .A2(_000_),
    .B(_105_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _363_ (.I(net157),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _364_ (.A1(net222),
    .A2(_074_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _365_ (.A1(_106_),
    .A2(_000_),
    .B(_107_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _366_ (.I0(net223),
    .I1(net158),
    .S(_073_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _367_ (.I(_108_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _368_ (.I(net159),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _369_ (.A1(net224),
    .A2(_074_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _370_ (.A1(_109_),
    .A2(_000_),
    .B(_110_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _371_ (.I0(net225),
    .I1(net160),
    .S(_073_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _372_ (.I(_111_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _373_ (.I0(net226),
    .I1(net161),
    .S(_073_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _374_ (.I(_112_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _375_ (.I0(net227),
    .I1(net162),
    .S(_073_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _376_ (.I(_113_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _377_ (.I(net163),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _378_ (.A1(net228),
    .A2(_074_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _379_ (.A1(_114_),
    .A2(_000_),
    .B(_115_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _380_ (.I(net165),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _381_ (.A1(net230),
    .A2(_074_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _382_ (.A1(_116_),
    .A2(_076_),
    .B(_117_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _383_ (.I(net166),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _384_ (.A1(net231),
    .A2(_074_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _385_ (.A1(_118_),
    .A2(_076_),
    .B(_119_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _386_ (.A1(net33),
    .A2(_069_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _387_ (.A1(net104),
    .A2(net99),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _388_ (.A1(net57),
    .A2(_069_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _389_ (.A1(net35),
    .A2(_069_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _390_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _391_ (.A1(net60),
    .A2(_069_),
    .B(_124_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _392_ (.I(_068_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _393_ (.A1(_066_),
    .A2(_126_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _394_ (.A1(net34),
    .A2(_069_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _395_ (.A1(_127_),
    .A2(_120_),
    .A3(_128_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _396_ (.A1(net41),
    .A2(_069_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _397_ (.A1(net52),
    .A2(_069_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _398_ (.A1(net44),
    .A2(_069_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _399_ (.A1(net62),
    .A2(_067_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _400_ (.A1(net59),
    .A2(_067_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _401_ (.A1(net63),
    .A2(_068_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _402_ (.A1(net58),
    .A2(net61),
    .B(_068_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _403_ (.A1(_133_),
    .A2(_134_),
    .A3(_135_),
    .A4(_136_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _404_ (.A1(_130_),
    .A2(_131_),
    .A3(_132_),
    .A4(_137_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _405_ (.A1(net46),
    .A2(_126_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _406_ (.A1(net43),
    .A2(_126_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _407_ (.A1(net42),
    .A2(_126_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _408_ (.A1(net45),
    .A2(_069_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _409_ (.A1(_139_),
    .A2(_140_),
    .A3(_141_),
    .A4(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _410_ (.A1(net53),
    .A2(_126_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _411_ (.A1(net54),
    .A2(_068_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _412_ (.A1(net55),
    .A2(_126_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _413_ (.A1(net38),
    .A2(_126_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _414_ (.A1(_144_),
    .A2(_145_),
    .A3(_146_),
    .A4(_147_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _415_ (.A1(net50),
    .A2(_126_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _416_ (.A1(net36),
    .A2(_068_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _417_ (.A1(net51),
    .A2(_068_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _418_ (.A1(net39),
    .A2(_126_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _419_ (.A1(_149_),
    .A2(_150_),
    .A3(_151_),
    .A4(_152_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _420_ (.A1(net37),
    .A2(net56),
    .B(_068_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _421_ (.A1(net48),
    .A2(_068_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _422_ (.A1(net47),
    .A2(net64),
    .B(_068_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _423_ (.A1(net40),
    .A2(net49),
    .B(_126_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _424_ (.A1(_154_),
    .A2(_155_),
    .A3(_156_),
    .A4(_157_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _425_ (.A1(_143_),
    .A2(_148_),
    .A3(_153_),
    .A4(_158_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _426_ (.A1(_125_),
    .A2(_129_),
    .A3(_138_),
    .A4(_159_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _427_ (.A1(_071_),
    .A2(_121_),
    .B(_160_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _428_ (.A1(net1),
    .A2(_120_),
    .B1(_161_),
    .B2(_075_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _429_ (.A1(net67),
    .A2(_076_),
    .A3(_121_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _430_ (.A1(_065_),
    .A2(_162_),
    .B(_163_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _431_ (.I(_065_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _432_ (.A1(net153),
    .A2(net142),
    .Z(_165_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _433_ (.A1(net78),
    .A2(_127_),
    .A3(_121_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _434_ (.A1(net2),
    .A2(_128_),
    .B1(_161_),
    .B2(_165_),
    .C(_166_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _435_ (.A1(_164_),
    .A2(_167_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _436_ (.A1(net153),
    .A2(net142),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _437_ (.A1(net164),
    .A2(_168_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _438_ (.A1(net3),
    .A2(_123_),
    .B1(_161_),
    .B2(_169_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _439_ (.A1(net89),
    .A2(_076_),
    .A3(_121_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _440_ (.A1(_065_),
    .A2(_170_),
    .B(_171_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _441_ (.A1(net164),
    .A2(net153),
    .A3(net142),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _442_ (.A1(net167),
    .A2(_172_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _443_ (.A1(net92),
    .A2(_127_),
    .A3(_121_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _444_ (.A1(net4),
    .A2(_150_),
    .B1(_161_),
    .B2(_173_),
    .C(_174_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _445_ (.A1(_164_),
    .A2(_175_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _446_ (.A1(net37),
    .A2(_070_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _447_ (.A1(net5),
    .A2(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _448_ (.A1(net167),
    .A2(net164),
    .A3(net153),
    .A4(net142),
    .Z(_178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _449_ (.A1(net168),
    .A2(_178_),
    .Z(_179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _450_ (.A1(_127_),
    .A2(_121_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _451_ (.A1(_161_),
    .A2(_179_),
    .B1(_180_),
    .B2(net93),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _452_ (.A1(_177_),
    .A2(_181_),
    .B(_164_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _453_ (.A1(net168),
    .A2(_178_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _454_ (.A1(net169),
    .A2(_182_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _455_ (.A1(net6),
    .A2(_147_),
    .B1(_161_),
    .B2(_183_),
    .C1(_180_),
    .C2(net94),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _456_ (.A1(_164_),
    .A2(_184_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _457_ (.A1(net7),
    .A2(_152_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _458_ (.A1(net169),
    .A2(net168),
    .A3(_178_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _459_ (.A1(net170),
    .A2(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _460_ (.A1(net95),
    .A2(_180_),
    .B1(_187_),
    .B2(_161_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _461_ (.A1(_185_),
    .A2(_188_),
    .B(_164_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _462_ (.A1(net40),
    .A2(_070_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _463_ (.A1(net170),
    .A2(net169),
    .A3(net168),
    .A4(_178_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _464_ (.A1(_085_),
    .A2(_190_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _465_ (.A1(net8),
    .A2(_189_),
    .B1(_161_),
    .B2(_191_),
    .C1(_180_),
    .C2(net96),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _466_ (.A1(_164_),
    .A2(_192_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _467_ (.I(_065_),
    .Z(_193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _468_ (.A1(net104),
    .A2(net100),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _469_ (.A1(_127_),
    .A2(_194_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _470_ (.A1(_160_),
    .A2(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _471_ (.A1(_085_),
    .A2(_190_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _472_ (.A1(net172),
    .A2(_197_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _473_ (.A1(_071_),
    .A2(_194_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _474_ (.A1(net9),
    .A2(_130_),
    .B1(_196_),
    .B2(_198_),
    .C1(_199_),
    .C2(net97),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _475_ (.A1(_193_),
    .A2(_200_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _476_ (.A1(net172),
    .A2(_197_),
    .B(net173),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _477_ (.A1(net173),
    .A2(net172),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _478_ (.A1(_085_),
    .A2(_190_),
    .A3(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _479_ (.A1(_201_),
    .A2(_203_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _480_ (.A1(_196_),
    .A2(_204_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _481_ (.A1(net10),
    .A2(_141_),
    .B1(_199_),
    .B2(net98),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _482_ (.A1(_205_),
    .A2(_206_),
    .B(_164_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _483_ (.A1(net143),
    .A2(_203_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _484_ (.A1(net11),
    .A2(_140_),
    .B1(_196_),
    .B2(_207_),
    .C1(_199_),
    .C2(net68),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _485_ (.A1(_193_),
    .A2(_208_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _486_ (.A1(_089_),
    .A2(_085_),
    .A3(_190_),
    .A4(_202_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _487_ (.A1(net144),
    .A2(_209_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _488_ (.A1(net12),
    .A2(_132_),
    .B1(_196_),
    .B2(_210_),
    .C1(_199_),
    .C2(net69),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _489_ (.A1(_193_),
    .A2(_211_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _490_ (.A1(net144),
    .A2(_209_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _491_ (.A1(net145),
    .A2(_212_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _492_ (.A1(net13),
    .A2(_142_),
    .B1(_196_),
    .B2(_213_),
    .C1(_199_),
    .C2(net70),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _493_ (.A1(_193_),
    .A2(_214_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _494_ (.A1(net145),
    .A2(_212_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _495_ (.A1(net146),
    .A2(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _496_ (.A1(net14),
    .A2(_139_),
    .B1(_196_),
    .B2(_216_),
    .C1(_199_),
    .C2(net71),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _497_ (.A1(_193_),
    .A2(_217_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _498_ (.A1(net146),
    .A2(net145),
    .A3(net144),
    .A4(_209_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _499_ (.A1(_094_),
    .A2(_218_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _500_ (.A1(_160_),
    .A2(_195_),
    .B1(_218_),
    .B2(_094_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _501_ (.I(net15),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _502_ (.A1(net47),
    .A2(_221_),
    .A3(_070_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _503_ (.A1(net72),
    .A2(_199_),
    .B1(_219_),
    .B2(_220_),
    .C(_222_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _504_ (.A1(_193_),
    .A2(_223_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _505_ (.A1(_096_),
    .A2(_219_),
    .Z(_224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _506_ (.A1(net16),
    .A2(_155_),
    .B1(_196_),
    .B2(_224_),
    .C1(_199_),
    .C2(net73),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _507_ (.A1(_193_),
    .A2(_225_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _508_ (.A1(net49),
    .A2(_070_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _509_ (.A1(net101),
    .A2(net104),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _510_ (.A1(_127_),
    .A2(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _511_ (.A1(_160_),
    .A2(_228_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _512_ (.A1(_096_),
    .A2(_219_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _513_ (.A1(net149),
    .A2(_230_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _514_ (.A1(_071_),
    .A2(_227_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _515_ (.A1(net17),
    .A2(_226_),
    .B1(_229_),
    .B2(_231_),
    .C1(_232_),
    .C2(net74),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _516_ (.A1(_193_),
    .A2(_233_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _517_ (.I(_229_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _518_ (.A1(net149),
    .A2(_230_),
    .B(net150),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _519_ (.A1(net149),
    .A2(net150),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _520_ (.A1(_096_),
    .A2(_094_),
    .A3(_218_),
    .A4(_236_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _521_ (.A1(_234_),
    .A2(_235_),
    .A3(_237_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _522_ (.A1(net18),
    .A2(_149_),
    .B1(_232_),
    .B2(net75),
    .C(_238_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _523_ (.A1(_193_),
    .A2(_239_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _524_ (.A1(net151),
    .A2(_237_),
    .Z(_240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _525_ (.A1(net19),
    .A2(_151_),
    .B1(_229_),
    .B2(_240_),
    .C1(_232_),
    .C2(net76),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _526_ (.A1(_193_),
    .A2(_241_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _527_ (.I(_065_),
    .Z(_242_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _528_ (.A1(net151),
    .A2(net152),
    .A3(_237_),
    .Z(_243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _529_ (.A1(net151),
    .A2(_237_),
    .B(net152),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _530_ (.A1(_234_),
    .A2(_243_),
    .A3(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _531_ (.A1(net20),
    .A2(_131_),
    .B1(_232_),
    .B2(net77),
    .C(_245_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _532_ (.A1(_242_),
    .A2(_246_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _533_ (.A1(net154),
    .A2(_243_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _534_ (.A1(net21),
    .A2(_144_),
    .B1(_229_),
    .B2(_247_),
    .C1(_232_),
    .C2(net79),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _535_ (.A1(_242_),
    .A2(_248_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _536_ (.A1(net154),
    .A2(_243_),
    .Z(_249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _537_ (.A1(net154),
    .A2(net155),
    .Z(_250_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _538_ (.A1(net151),
    .A2(net152),
    .A3(_237_),
    .A4(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _539_ (.A1(net155),
    .A2(_249_),
    .B(_251_),
    .C(_229_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _540_ (.A1(net22),
    .A2(_145_),
    .B1(_232_),
    .B2(net80),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _541_ (.A1(_252_),
    .A2(_253_),
    .B(_164_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _542_ (.A1(_104_),
    .A2(_251_),
    .Z(_254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _543_ (.A1(net23),
    .A2(_146_),
    .B1(_229_),
    .B2(_254_),
    .C1(_232_),
    .C2(net81),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _544_ (.A1(_242_),
    .A2(_255_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _545_ (.A1(net56),
    .A2(_070_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _546_ (.A1(_104_),
    .A2(_251_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _547_ (.A1(net157),
    .A2(_257_),
    .Z(_258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _548_ (.A1(net24),
    .A2(_256_),
    .B1(_229_),
    .B2(_258_),
    .C1(_232_),
    .C2(net82),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _549_ (.A1(_242_),
    .A2(_259_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _550_ (.A1(net104),
    .A2(net102),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _551_ (.A1(_127_),
    .A2(_260_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _552_ (.A1(_160_),
    .A2(_261_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _553_ (.A1(net157),
    .A2(_257_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _554_ (.A1(net158),
    .A2(_263_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _555_ (.A1(_071_),
    .A2(_260_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _556_ (.A1(net25),
    .A2(_122_),
    .B1(_262_),
    .B2(_264_),
    .C1(_265_),
    .C2(net83),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _557_ (.A1(_242_),
    .A2(_266_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _558_ (.A1(net58),
    .A2(_070_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _559_ (.A1(net157),
    .A2(net158),
    .A3(_257_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _560_ (.I(_262_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _561_ (.A1(net158),
    .A2(net159),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _562_ (.A1(_104_),
    .A2(_106_),
    .A3(_251_),
    .A4(_270_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _563_ (.A1(_109_),
    .A2(_268_),
    .B(_269_),
    .C(_271_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _564_ (.A1(net26),
    .A2(_267_),
    .B1(_265_),
    .B2(net84),
    .C(_272_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _565_ (.A1(_242_),
    .A2(_273_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _566_ (.A1(net160),
    .A2(_271_),
    .Z(_274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _567_ (.A1(net27),
    .A2(_134_),
    .B1(_262_),
    .B2(_274_),
    .C1(_265_),
    .C2(net85),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _568_ (.A1(_242_),
    .A2(_275_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _569_ (.A1(net160),
    .A2(net161),
    .A3(_271_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _570_ (.A1(net160),
    .A2(_271_),
    .B(net161),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _571_ (.A1(_269_),
    .A2(_277_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _572_ (.I(net28),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _573_ (.A1(net60),
    .A2(_279_),
    .A3(_070_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _574_ (.A1(net86),
    .A2(_265_),
    .B1(_276_),
    .B2(_278_),
    .C(_280_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _575_ (.A1(_242_),
    .A2(_281_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _576_ (.A1(net61),
    .A2(_070_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _577_ (.A1(net162),
    .A2(_276_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _578_ (.A1(net29),
    .A2(_282_),
    .B1(_262_),
    .B2(_283_),
    .C1(_265_),
    .C2(net87),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _579_ (.A1(_242_),
    .A2(_284_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _580_ (.A1(net160),
    .A2(net161),
    .A3(net162),
    .A4(_271_),
    .Z(_285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _581_ (.A1(net163),
    .A2(_285_),
    .Z(_286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _582_ (.A1(net30),
    .A2(_133_),
    .B1(_262_),
    .B2(_286_),
    .C1(_265_),
    .C2(net88),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _583_ (.A1(_242_),
    .A2(_287_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _584_ (.A1(net163),
    .A2(net165),
    .A3(_285_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _585_ (.A1(net160),
    .A2(net161),
    .A3(net162),
    .A4(_271_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _586_ (.A1(_114_),
    .A2(_289_),
    .B(_116_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _587_ (.A1(_262_),
    .A2(_288_),
    .A3(_290_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _588_ (.A1(net31),
    .A2(_135_),
    .B1(_265_),
    .B2(net90),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _589_ (.A1(_291_),
    .A2(_292_),
    .B(_164_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _590_ (.A1(net163),
    .A2(net165),
    .A3(net166),
    .A4(_285_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _591_ (.A1(_114_),
    .A2(_116_),
    .A3(_289_),
    .B(_118_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _592_ (.A1(_262_),
    .A2(_293_),
    .A3(_294_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _593_ (.A1(net64),
    .A2(_070_),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _594_ (.A1(net32),
    .A2(_296_),
    .B1(_265_),
    .B2(net91),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _595_ (.A1(_295_),
    .A2(_297_),
    .B(_164_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _596_ (.D(_000_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net206));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _597_ (.D(_001_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net207));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _598_ (.D(_002_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net218));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _599_ (.D(_003_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _600_ (.D(_004_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _601_ (.D(_005_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net233));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _602_ (.D(_006_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net234));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _603_ (.D(_007_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net235));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _604_ (.D(_008_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net236));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _605_ (.D(_009_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net237));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _606_ (.D(_010_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net238));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _607_ (.D(_011_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net208));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _608_ (.D(_012_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net209));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _609_ (.D(_013_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net210));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _610_ (.D(_014_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net211));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _611_ (.D(_015_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net212));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _612_ (.D(_016_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net213));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _613_ (.D(_017_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net214));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _614_ (.D(_018_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net215));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _615_ (.D(_019_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net216));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _616_ (.D(_020_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net217));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _617_ (.D(_021_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net219));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _618_ (.D(_022_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net220));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _619_ (.D(_023_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net221));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _620_ (.D(_024_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net222));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _621_ (.D(_025_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net223));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _622_ (.D(_026_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _623_ (.D(_027_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _624_ (.D(_028_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _625_ (.D(_029_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _626_ (.D(_030_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _627_ (.D(_031_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net230));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _628_ (.D(_032_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net231));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _629_ (.D(_033_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _630_ (.D(_034_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _631_ (.D(_035_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net164));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _632_ (.D(_036_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net167));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _633_ (.D(_037_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net168));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _634_ (.D(_038_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(net169));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _635_ (.D(_039_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net170));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _636_ (.D(_040_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net171));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _637_ (.D(_041_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net172));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _638_ (.D(_042_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net173));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _639_ (.D(_043_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _640_ (.D(_044_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _641_ (.D(_045_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _642_ (.D(_046_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _643_ (.D(_047_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net147));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _644_ (.D(_048_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _645_ (.D(_049_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net149));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _646_ (.D(_050_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _647_ (.D(_051_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _648_ (.D(_052_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net152));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _649_ (.D(_053_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net154));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _650_ (.D(_054_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net155));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _651_ (.D(_055_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net156));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _652_ (.D(_056_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net157));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _653_ (.D(_057_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net158));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _654_ (.D(_058_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _655_ (.D(_059_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net160));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _656_ (.D(_060_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _657_ (.D(_061_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net162));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _658_ (.D(_062_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net163));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _659_ (.D(_063_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net165));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _660_ (.D(_064_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _703_ (.I(net239),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _704_ (.I(net241),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _705_ (.I(net242),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _706_ (.I(net242),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _707_ (.I(net239),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _708_ (.I(net243),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _709_ (.I(net240),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _710_ (.I(net241),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _711_ (.I(net242),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _712_ (.I(net242),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _713_ (.I(net239),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _714_ (.I(net239),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _715_ (.I(net239),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _716_ (.I(net241),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _717_ (.I(net241),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _718_ (.I(net243),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _719_ (.I(net239),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _720_ (.I(net239),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _721_ (.I(net239),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _722_ (.I(net240),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _723_ (.I(net241),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _724_ (.I(net240),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _725_ (.I(net241),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _726_ (.I(net240),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _727_ (.I(net241),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _728_ (.I(net240),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _729_ (.I(net241),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _730_ (.I(net239),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _731_ (.I(net239),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _732_ (.I(net240),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _733_ (.I(net240),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _734_ (.I(net243),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _735_ (.I(net241),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _736_ (.I(net240),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _737_ (.I(net240),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _738_ (.I(net243),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _739_ (.I(net241),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _740_ (.I(net142),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _741_ (.I(net153),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _742_ (.I(net164),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _743_ (.I(net167),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _744_ (.I(net168),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _745_ (.I(net169),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _746_ (.I(net170),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _747_ (.I(net171),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _748_ (.I(net172),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _749_ (.I(net173),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _750_ (.I(net143),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _751_ (.I(net144),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _752_ (.I(net145),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _753_ (.I(net146),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _754_ (.I(net147),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _755_ (.I(net148),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _756_ (.I(net149),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _757_ (.I(net150),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _758_ (.I(net151),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _759_ (.I(net152),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _760_ (.I(net154),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _761_ (.I(net155),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _762_ (.I(net156),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _763_ (.I(net157),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _764_ (.I(net158),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _765_ (.I(net159),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _766_ (.I(net160),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _767_ (.I(net161),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _768_ (.I(net162),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _769_ (.I(net163),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _770_ (.I(net165),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _771_ (.I(net166),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(la_data_in[32]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(la_data_in[33]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(la_data_in[34]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(la_data_in[35]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(la_data_in[36]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(la_data_in[37]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(la_data_in[38]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(la_data_in[39]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(la_data_in[40]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(la_data_in[41]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(la_data_in[42]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(la_data_in[43]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(la_data_in[44]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(la_data_in[45]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(la_data_in[46]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(la_data_in[47]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(la_data_in[48]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(la_data_in[49]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(la_data_in[50]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(la_data_in[51]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(la_data_in[52]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(la_data_in[53]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(la_data_in[54]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(la_data_in[55]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(la_data_in[56]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(la_data_in[57]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(la_data_in[58]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(la_data_in[59]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(la_data_in[60]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(la_data_in[61]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(la_data_in[62]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(la_data_in[63]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(la_oenb[32]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(la_oenb[33]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(la_oenb[34]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(la_oenb[35]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(la_oenb[36]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(la_oenb[37]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(la_oenb[38]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input40 (.I(la_oenb[39]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(la_oenb[40]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(la_oenb[41]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(la_oenb[42]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(la_oenb[43]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input45 (.I(la_oenb[44]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input46 (.I(la_oenb[45]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input47 (.I(la_oenb[46]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input48 (.I(la_oenb[47]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input49 (.I(la_oenb[48]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input50 (.I(la_oenb[49]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(la_oenb[50]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input52 (.I(la_oenb[51]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(la_oenb[52]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input54 (.I(la_oenb[53]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input55 (.I(la_oenb[54]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input56 (.I(la_oenb[55]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input57 (.I(la_oenb[56]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(la_oenb[57]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input59 (.I(la_oenb[58]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(la_oenb[59]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input61 (.I(la_oenb[60]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input62 (.I(la_oenb[61]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input63 (.I(la_oenb[62]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input64 (.I(la_oenb[63]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(wb_rst_i),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(wbs_cyc_i),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input67 (.I(wbs_dat_i[0]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(wbs_dat_i[10]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(wbs_dat_i[11]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(wbs_dat_i[12]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input71 (.I(wbs_dat_i[13]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(wbs_dat_i[14]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input73 (.I(wbs_dat_i[15]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(wbs_dat_i[16]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input75 (.I(wbs_dat_i[17]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input76 (.I(wbs_dat_i[18]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input77 (.I(wbs_dat_i[19]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input78 (.I(wbs_dat_i[1]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input79 (.I(wbs_dat_i[20]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(wbs_dat_i[21]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input81 (.I(wbs_dat_i[22]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input82 (.I(wbs_dat_i[23]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input83 (.I(wbs_dat_i[24]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input84 (.I(wbs_dat_i[25]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input85 (.I(wbs_dat_i[26]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input86 (.I(wbs_dat_i[27]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input87 (.I(wbs_dat_i[28]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input88 (.I(wbs_dat_i[29]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input89 (.I(wbs_dat_i[2]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(wbs_dat_i[30]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input91 (.I(wbs_dat_i[31]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input92 (.I(wbs_dat_i[3]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input93 (.I(wbs_dat_i[4]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input94 (.I(wbs_dat_i[5]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(wbs_dat_i[6]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input96 (.I(wbs_dat_i[7]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input97 (.I(wbs_dat_i[8]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input98 (.I(wbs_dat_i[9]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(wbs_sel_i[0]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input100 (.I(wbs_sel_i[1]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(wbs_sel_i[2]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(wbs_sel_i[3]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input103 (.I(wbs_stb_i),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input104 (.I(wbs_we_i),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output105 (.I(net105),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output106 (.I(net106),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output107 (.I(net107),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output108 (.I(net108),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output109 (.I(net109),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output110 (.I(net110),
    .Z(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output111 (.I(net111),
    .Z(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output112 (.I(net112),
    .Z(io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output113 (.I(net113),
    .Z(io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output114 (.I(net114),
    .Z(io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output115 (.I(net115),
    .Z(io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output116 (.I(net116),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output117 (.I(net117),
    .Z(io_oeb[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output118 (.I(net118),
    .Z(io_oeb[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output119 (.I(net119),
    .Z(io_oeb[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output120 (.I(net120),
    .Z(io_oeb[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output121 (.I(net121),
    .Z(io_oeb[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output122 (.I(net122),
    .Z(io_oeb[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output123 (.I(net123),
    .Z(io_oeb[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output124 (.I(net124),
    .Z(io_oeb[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output125 (.I(net125),
    .Z(io_oeb[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output126 (.I(net126),
    .Z(io_oeb[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(io_oeb[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(io_oeb[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(io_oeb[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output131 (.I(net131),
    .Z(io_oeb[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output132 (.I(net132),
    .Z(io_oeb[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(io_oeb[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(io_oeb[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net159),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net186),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output192 (.I(net192),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output193 (.I(net193),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output194 (.I(net194),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output195 (.I(net195),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output196 (.I(net196),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output197 (.I(net197),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output198 (.I(net198),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output199 (.I(net199),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output200 (.I(net200),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output201 (.I(net201),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output202 (.I(net202),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output203 (.I(net203),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output204 (.I(net204),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output205 (.I(net205),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output206 (.I(net206),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output207 (.I(net207),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output208 (.I(net208),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output209 (.I(net209),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output210 (.I(net210),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output211 (.I(net211),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output212 (.I(net212),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output213 (.I(net213),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output214 (.I(net214),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output215 (.I(net215),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output216 (.I(net216),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output217 (.I(net217),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output218 (.I(net218),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output219 (.I(net219),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output220 (.I(net220),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output221 (.I(net221),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output222 (.I(net222),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output223 (.I(net223),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output224 (.I(net224),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output225 (.I(net225),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output226 (.I(net226),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output227 (.I(net227),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output228 (.I(net228),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output229 (.I(net229),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output230 (.I(net230),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output231 (.I(net231),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output232 (.I(net232),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output233 (.I(net233),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output234 (.I(net234),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output235 (.I(net235),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output236 (.I(net236),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output237 (.I(net237),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output238 (.I(net238),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout239 (.I(net240),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout240 (.I(net65),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout241 (.I(net242),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout242 (.I(net243),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout243 (.I(net65),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__596__D (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A2 (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__A2 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A2 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__B (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__B (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__B (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__I (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__I (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__I (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__593__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__576__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__A3 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__558__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A3 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__S (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__I (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__I (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__S (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__S (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__S (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__S (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__B2 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A1 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__S (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__486__A2 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__A2 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__B2 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__A1 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__A1 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__591__A2 (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__586__B (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__A1 (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__A1 (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__B (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__A2 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A2 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__A2 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__A2 (.I(_132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A3 (.I(_132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__A2 (.I(_133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A1 (.I(_133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A2 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A2 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A2 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A3 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__A2 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__A1 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__A2 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__A2 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__A2 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__A4 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__A2 (.I(_144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A1 (.I(_144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__A2 (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A2 (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__A2 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A3 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A2 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A2 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A2 (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A4 (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__552__A1 (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A1 (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__A1 (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__A1 (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__B (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__B2 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__B1 (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__595__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A1 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__A1 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__B (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A1 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__A1 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__A1 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__C1 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A2 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__C1 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__B1 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__486__A3 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__A2 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__A2 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A2 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__B1 (.I(_196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A2 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__B1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__C1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A4 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__A2 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__A2 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__A3 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__B1 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__A2 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__B1 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__B1 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__C (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__B1 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__B1 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__I (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__B1 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__C1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__C1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__C1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__B1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__C1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__B1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__C1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__A3 (.I(_237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A2 (.I(_237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A3 (.I(_237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__A2 (.I(_237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__A3 (.I(_237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__579__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__565__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__549__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__A2 (.I(_243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__A2 (.I(_243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__A2 (.I(_243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A3 (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A2 (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__A2 (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__B (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__A2 (.I(_253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A3 (.I(_257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__A2 (.I(_257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__547__A2 (.I(_257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__592__A1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__A1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__B1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__B1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__B1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__I (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__B1 (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__B1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__B1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__C1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__C1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__A2 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__C1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__C1 (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A4 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A4 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__A2 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__A3 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__A2 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__C (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__C (.I(_280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(la_data_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(la_data_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(la_data_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(la_data_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(la_data_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(la_data_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(la_data_in[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(la_data_in[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(la_data_in[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(la_data_in[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(la_data_in[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(la_data_in[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(la_data_in[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(la_data_in[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(la_data_in[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(la_data_in[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(la_data_in[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(la_data_in[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(la_data_in[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(la_data_in[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_data_in[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_data_in[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(la_data_in[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(la_data_in[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(la_data_in[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(la_data_in[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(la_data_in[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(la_data_in[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(la_data_in[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(la_data_in[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(la_data_in[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(la_oenb[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(la_oenb[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_oenb[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(la_oenb[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(la_oenb[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(la_oenb[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(la_oenb[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(la_oenb[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(la_oenb[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(la_oenb[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(la_oenb[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(la_oenb[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(la_oenb[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(la_oenb[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(la_oenb[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(la_oenb[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(la_oenb[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(la_oenb[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(la_oenb[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(la_oenb[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(la_oenb[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(la_oenb[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(la_oenb[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(la_oenb[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(la_oenb[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(la_oenb[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(la_oenb[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(la_oenb[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(la_oenb[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(la_oenb[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(la_oenb[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(la_oenb[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(wbs_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(wbs_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(wbs_sel_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(wbs_sel_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A2 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__558__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__576__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__593__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout243_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__C2 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__C2 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__C2 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__C2 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__C2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__C2 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__B2 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__C2 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__B2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__C2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__C2 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__C2 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__C2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__C2 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__C2 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__C2 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__B2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__B2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__B2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__C2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__C2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__C2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__B2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__A2 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A2 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__A2 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__740__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A4 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A3 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__750__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A3 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__I1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__752__I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A2 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__I1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__753__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A1 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A1 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__I1 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__754__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__755__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__756__I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__757__I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__A2 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__B (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__I1 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__758__I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__I1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__759__I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__B (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__741__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A3 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__I1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__760__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__A1 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__A1 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__A1 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__I1 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__761__I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__A1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__762__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__763__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__547__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__764__I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A2 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__I1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__765__I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__766__I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__I1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__767__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__B (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__I1 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__768__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A3 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A3 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__577__A1 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__I1 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__769__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__742__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A2 (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A1 (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__A1 (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__I1 (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__A2 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__A2 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__771__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__A3 (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__I1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__744__I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A3 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__A1 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A1 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__I1 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__745__I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A1 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A1 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__I1 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A1 (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A1 (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__I1 (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__747__I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__748__I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__A2 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__I1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__749__I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__B (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__I1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__I0 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__I0 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__I0 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A1 (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I0 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__I0 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__I0 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I0 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__I0 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__I0 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I0 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A1 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__I0 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__I0 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__I0 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__I0 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A1 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A1 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output231_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A1 (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output232_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__I0 (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output233_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__I0 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output234_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__I0 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output235_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__I0 (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A1 (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__I0 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output238_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__I0 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__731__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__721__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__720__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__715__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__703__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__730__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__719__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__714__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout239_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__736__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__733__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__728__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__726__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__724__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__722__I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__739__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__735__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__727__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__725__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__723__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__717__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__704__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__706__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__711__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__712__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout241_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__705__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__738__I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__718__I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__708__I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout242_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__601__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__602__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__613__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__616__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__625__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__634__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__598__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__599__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__615__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__635__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__614__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__620__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__621__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__622__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__630__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__649__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__650__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__651__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__654__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__596__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__604__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__633__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__653__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__617__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__618__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__619__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__640__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__643__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__648__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__655__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__597__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__629__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__631__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__645__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__652__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__607__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__612__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__624__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__627__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__636__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__637__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__638__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__639__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__641__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__642__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__644__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__660__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__603__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__605__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__606__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__609__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__610__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__611__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__626__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__658__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__659__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 assign io_oeb[37] = net244;
 assign io_out[32] = net245;
 assign io_out[33] = net246;
 assign io_out[34] = net247;
 assign io_out[35] = net248;
 assign io_out[36] = net249;
 assign io_out[37] = net250;
 assign irq[0] = net251;
 assign irq[1] = net252;
 assign irq[2] = net253;
 assign la_data_out[32] = net254;
 assign la_data_out[33] = net255;
 assign la_data_out[34] = net256;
 assign la_data_out[35] = net257;
 assign la_data_out[36] = net258;
 assign la_data_out[37] = net259;
 assign la_data_out[38] = net260;
 assign la_data_out[39] = net261;
 assign la_data_out[40] = net262;
 assign la_data_out[41] = net263;
 assign la_data_out[42] = net264;
 assign la_data_out[43] = net265;
 assign la_data_out[44] = net266;
 assign la_data_out[45] = net267;
 assign la_data_out[46] = net268;
 assign la_data_out[47] = net269;
 assign la_data_out[48] = net270;
 assign la_data_out[49] = net271;
 assign la_data_out[50] = net272;
 assign la_data_out[51] = net273;
 assign la_data_out[52] = net274;
 assign la_data_out[53] = net275;
 assign la_data_out[54] = net276;
 assign la_data_out[55] = net277;
 assign la_data_out[56] = net278;
 assign la_data_out[57] = net279;
 assign la_data_out[58] = net280;
 assign la_data_out[59] = net281;
 assign la_data_out[60] = net282;
 assign la_data_out[61] = net283;
 assign la_data_out[62] = net284;
 assign la_data_out[63] = net285;
endmodule

