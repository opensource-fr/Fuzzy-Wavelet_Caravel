VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.040 4.000 209.160 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.240 4.000 276.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.360 4.000 249.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.640 596.000 578.760 599.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 211.400 4.000 212.520 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.000 596.000 330.120 599.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 113.960 599.000 115.080 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.080 1.000 172.200 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 596.000 135.240 599.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 265.160 4.000 266.280 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 597.800 599.000 598.920 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.200 596.000 481.320 599.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.800 596.000 346.920 599.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.560 596.000 568.680 599.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 596.000 10.920 599.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 1.000 81.480 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 596.000 74.760 599.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 596.000 98.280 599.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 63.560 599.000 64.680 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.200 4.000 145.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.240 596.000 24.360 599.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 584.360 599.000 585.480 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.200 4.000 61.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.720 1.000 420.840 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.080 596.000 88.200 599.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.880 1.000 357.000 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 587.720 4.000 588.840 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.320 596.000 538.440 599.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.400 596.000 128.520 599.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.280 4.000 155.400 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 97.160 599.000 98.280 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 251.720 4.000 252.840 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.320 1.000 538.440 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.360 4.000 585.480 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.480 4.000 138.600 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 157.640 599.000 158.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.360 1.000 585.480 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.440 596.000 511.560 599.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.520 596.000 17.640 599.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 409.640 4.000 410.760 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 376.040 4.000 377.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 449.960 4.000 451.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.800 1.000 514.920 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 587.720 1.000 588.840 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.920 596.000 320.040 599.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 345.800 4.000 346.920 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 596.000 57.960 599.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.480 4.000 474.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.640 1.000 242.760 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 46.760 599.000 47.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.080 1.000 508.200 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 1.000 57.960 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 150.920 599.000 152.040 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 56.840 4.000 57.960 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 134.120 599.000 135.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.400 1.000 212.520 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.000 1.000 498.120 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.560 4.000 400.680 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 560.840 4.000 561.960 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 596.000 121.800 599.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.120 1.000 387.240 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 19.880 4.000 21.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 416.360 599.000 417.480 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 93.800 599.000 94.920 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.280 4.000 491.400 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.560 4.000 232.680 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.720 596.000 336.840 599.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.840 1.000 561.960 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 503.720 4.000 504.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 201.320 599.000 202.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 596.000 0.840 599.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 577.640 599.000 578.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 596.000 289.800 599.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 33.320 599.000 34.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 241.640 599.000 242.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 238.280 599.000 239.400 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 113.960 4.000 115.080 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.360 596.000 585.480 599.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 527.240 599.000 528.360 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 591.080 599.000 592.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 443.240 4.000 444.360 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.920 1.000 236.040 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 497.000 599.000 498.120 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 1.000 68.040 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.720 1.000 504.840 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.840 1.000 393.960 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 1.000 41.160 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.640 1.000 410.760 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.880 1.000 273.000 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.320 1.000 202.440 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.360 4.000 81.480 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.880 596.000 441.000 599.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 596.000 279.720 599.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.720 1.000 252.840 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.080 596.000 424.200 599.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.240 1.000 444.360 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.760 596.000 383.880 599.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.560 1.000 568.680 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 550.760 596.000 551.880 599.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 127.400 599.000 128.520 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.720 596.000 504.840 599.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 191.240 599.000 192.360 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.560 1.000 400.680 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 389.480 599.000 390.600 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 1.000 145.320 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 560.840 599.000 561.960 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 557.480 599.000 558.600 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 429.800 599.000 430.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.520 4.000 17.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.600 4.000 27.720 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 339.080 4.000 340.200 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.040 596.000 377.160 599.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 1.000 155.400 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 305.480 4.000 306.600 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 419.720 4.000 420.840 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.640 4.000 242.760 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 1.000 185.640 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.640 596.000 242.760 599.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.840 596.000 561.960 599.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.960 1.000 283.080 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.600 4.000 363.720 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 87.080 599.000 88.200 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 218.120 599.000 219.240 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 416.360 4.000 417.480 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 596.000 138.600 599.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 120.680 599.000 121.800 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 453.320 599.000 454.440 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 265.160 599.000 266.280 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.680 596.000 457.800 599.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.480 596.000 306.600 599.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.160 4.000 98.280 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.320 596.000 370.440 599.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.040 4.000 545.160 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.800 596.000 262.920 599.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 144.200 599.000 145.320 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.600 1.000 195.720 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.400 4.000 44.520 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.120 4.000 219.240 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 456.680 4.000 457.800 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 402.920 4.000 404.040 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.760 596.000 47.880 599.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 530.600 4.000 531.720 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.120 596.000 303.240 599.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 510.440 599.000 511.560 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 596.000 185.640 599.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 596.000 249.480 599.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 325.640 599.000 326.760 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 1.000 209.160 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 1.000 289.800 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.320 4.000 202.440 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 369.320 599.000 370.440 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 6.440 599.000 7.560 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 567.560 4.000 568.680 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 433.160 599.000 434.280 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.320 1.000 370.440 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.960 596.000 283.080 599.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 596.000 81.480 599.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 596.000 51.240 599.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 596.000 239.400 599.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.240 1.000 276.360 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 312.200 4.000 313.320 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.640 596.000 494.760 599.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.520 4.000 185.640 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.000 4.000 162.120 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 177.800 4.000 178.920 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 16.520 599.000 17.640 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 1.000 219.240 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 544.040 599.000 545.160 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 1.000 105.000 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.640 596.000 158.760 599.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.840 596.000 225.960 599.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.520 1.000 353.640 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 3.080 4.000 4.200 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 1.000 121.800 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 214.760 599.000 215.880 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 596.000 178.920 599.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.040 596.000 545.160 599.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.520 596.000 521.640 599.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 318.920 599.000 320.040 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.440 1.000 427.560 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 433.160 4.000 434.280 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.720 596.000 168.840 599.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 248.360 599.000 249.480 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 513.800 4.000 514.920 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 329.000 599.000 330.120 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.400 596.000 296.520 599.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.160 596.000 266.280 599.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.560 1.000 316.680 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 278.600 599.000 279.720 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.080 596.000 592.200 599.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 594.440 4.000 595.560 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 376.040 599.000 377.160 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 1.000 178.920 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 174.440 599.000 175.560 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 103.880 4.000 105.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 73.640 599.000 74.760 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.960 596.000 367.080 599.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 473.480 599.000 474.600 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.440 1.000 259.560 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 466.760 4.000 467.880 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 271.880 599.000 273.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 224.840 4.000 225.960 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.520 596.000 353.640 599.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 110.600 599.000 111.720 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.040 1.000 293.160 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.640 596.000 326.760 599.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 480.200 599.000 481.320 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 231.560 599.000 232.680 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 9.800 599.000 10.920 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 80.360 599.000 81.480 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.320 4.000 34.440 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.320 4.000 538.440 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 271.880 4.000 273.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 503.720 599.000 504.840 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 1.000 34.440 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 1.000 249.480 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.800 596.000 94.920 599.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.400 1.000 548.520 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.440 4.000 427.560 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 1.000 138.600 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.040 1.000 545.160 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.440 596.000 343.560 599.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 596.000 209.160 599.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.640 4.000 578.760 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.160 596.000 434.280 599.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 9.800 4.000 10.920 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.120 596.000 471.240 599.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.080 596.000 256.200 599.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 83.720 4.000 84.840 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 352.520 599.000 353.640 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 409.640 599.000 410.760 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 533.960 599.000 535.080 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 547.400 4.000 548.520 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.920 596.000 488.040 599.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.000 1.000 162.120 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.520 1.000 521.640 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 40.040 599.000 41.160 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.440 4.000 91.560 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.760 596.000 215.880 599.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.040 1.000 377.160 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 281.960 599.000 283.080 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 224.840 599.000 225.960 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 423.080 599.000 424.200 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 335.720 599.000 336.840 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 596.000 232.680 599.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.200 4.000 481.320 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.880 1.000 441.000 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.240 1.000 528.360 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.720 1.000 84.840 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.640 4.000 74.760 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 596.000 41.160 599.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 50.120 599.000 51.240 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 596.000 115.080 599.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.240 4.000 528.360 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.240 596.000 528.360 599.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.600 596.000 447.720 599.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.720 1.000 168.840 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 335.720 4.000 336.840 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.600 1.000 531.720 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 322.280 4.000 323.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.240 1.000 108.360 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 369.320 4.000 370.440 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 567.560 599.000 568.680 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 597.800 596.000 598.920 599.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 513.800 599.000 514.920 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 493.640 599.000 494.760 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 486.920 599.000 488.040 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.480 1.000 306.600 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 596.000 105.000 599.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.520 1.000 17.640 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.080 1.000 4.200 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.440 596.000 7.560 599.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.200 1.000 313.320 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.440 4.000 259.560 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.000 4.000 330.120 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.080 4.000 172.200 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 596.000 219.240 599.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 379.400 4.000 380.520 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 1.000 115.080 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.160 1.000 266.280 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 298.760 4.000 299.880 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.200 1.000 481.320 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.840 1.000 225.960 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 439.880 4.000 441.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 288.680 599.000 289.800 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 399.560 599.000 400.680 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.400 1.000 464.520 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.960 596.000 199.080 599.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.440 1.000 595.560 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 382.760 599.000 383.880 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.280 596.000 407.400 599.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 305.480 599.000 306.600 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.680 1.000 457.800 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 533.960 596.000 535.080 599.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 56.840 599.000 57.960 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.240 596.000 360.360 599.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.120 1.000 555.240 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.040 4.000 293.160 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 1.000 74.760 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 302.120 599.000 303.240 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 570.920 4.000 572.040 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 392.840 599.000 393.960 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.560 1.000 148.680 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.920 1.000 572.040 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.240 4.000 108.360 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.800 596.000 514.920 599.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 456.680 599.000 457.800 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.920 596.000 152.040 599.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.120 4.000 387.240 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 103.880 599.000 105.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.600 596.000 111.720 599.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 208.040 599.000 209.160 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.560 596.000 400.680 599.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.880 596.000 273.000 599.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 596.000 34.440 599.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 1.000 51.240 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.720 1.000 336.840 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 439.880 599.000 441.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 406.280 599.000 407.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.400 1.000 380.520 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 359.240 599.000 360.360 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 184.520 599.000 185.640 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.640 1.000 578.760 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.040 4.000 41.160 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 352.520 4.000 353.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.080 1.000 340.200 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.560 1.000 484.680 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 137.480 599.000 138.600 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 596.000 71.400 599.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.000 1.000 330.120 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 1.000 61.320 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.320 596.000 202.440 599.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 345.800 599.000 346.920 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 574.280 599.000 575.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 66.920 4.000 68.040 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 234.920 4.000 236.040 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 255.080 599.000 256.200 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.760 1.000 467.880 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.400 596.000 464.520 599.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.960 1.000 451.080 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.680 4.000 289.800 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 1.000 27.720 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 -0.280 599.000 0.840 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 161.000 599.000 162.120 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 596.000 192.360 599.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 520.520 599.000 521.640 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 463.400 4.000 464.520 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.080 4.000 508.200 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.560 4.000 484.680 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 1.000 21.000 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.040 4.000 125.160 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 312.200 599.000 313.320 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.800 1.000 346.920 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.640 596.000 410.760 599.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.480 596.000 558.600 599.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.960 596.000 31.080 599.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 1.000 91.560 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.560 4.000 148.680 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.280 596.000 575.400 599.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 355.880 4.000 357.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 470.120 599.000 471.240 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 197.960 599.000 199.080 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.360 1.000 417.480 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.000 596.000 498.120 599.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 596.000 145.320 599.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.880 1.000 189.000 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 365.960 599.000 367.080 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.280 1.000 491.400 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 177.800 599.000 178.920 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.560 4.000 316.680 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 23.240 599.000 24.360 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 1.000 98.280 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.760 1.000 299.880 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 261.800 599.000 262.920 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.480 596.000 474.600 599.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 537.320 599.000 538.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 29.960 599.000 31.080 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.680 4.000 121.800 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 342.440 599.000 343.560 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 1.000 10.920 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 550.760 599.000 551.880 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.320 596.000 454.440 599.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 70.280 599.000 71.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 429.800 596.000 430.920 599.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 167.720 4.000 168.840 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 187.880 4.000 189.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.920 1.000 404.040 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 1.000 0.840 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.480 1.000 474.600 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 281.960 4.000 283.080 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.520 4.000 521.640 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.000 596.000 162.120 599.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.600 4.000 195.720 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.040 1.000 125.160 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.400 1.000 44.520 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.200 596.000 313.320 599.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 596.000 175.560 599.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.280 1.000 323.400 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.360 596.000 417.480 599.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 167.720 599.000 168.840 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 392.840 4.000 393.960 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 463.400 599.000 464.520 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.760 1.000 131.880 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 1.000 232.680 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.120 4.000 51.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 446.600 599.000 447.720 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.600 1.000 363.720 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.840 596.000 393.960 599.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.480 596.000 390.600 599.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 554.120 4.000 555.240 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.560 596.000 64.680 599.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.160 1.000 434.280 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 130.760 4.000 131.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.000 4.000 498.120 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 295.400 599.000 296.520 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 593.040 585.610 ;
      LAYER Metal2 ;
        RECT 1.140 595.700 6.140 596.820 ;
        RECT 7.860 595.700 9.500 596.820 ;
        RECT 11.220 595.700 16.220 596.820 ;
        RECT 17.940 595.700 22.940 596.820 ;
        RECT 24.660 595.700 29.660 596.820 ;
        RECT 31.380 595.700 33.020 596.820 ;
        RECT 34.740 595.700 39.740 596.820 ;
        RECT 41.460 595.700 46.460 596.820 ;
        RECT 48.180 595.700 49.820 596.820 ;
        RECT 51.540 595.700 56.540 596.820 ;
        RECT 58.260 595.700 63.260 596.820 ;
        RECT 64.980 595.700 69.980 596.820 ;
        RECT 71.700 595.700 73.340 596.820 ;
        RECT 75.060 595.700 80.060 596.820 ;
        RECT 81.780 595.700 86.780 596.820 ;
        RECT 88.500 595.700 93.500 596.820 ;
        RECT 95.220 595.700 96.860 596.820 ;
        RECT 98.580 595.700 103.580 596.820 ;
        RECT 105.300 595.700 110.300 596.820 ;
        RECT 112.020 595.700 113.660 596.820 ;
        RECT 115.380 595.700 120.380 596.820 ;
        RECT 122.100 595.700 127.100 596.820 ;
        RECT 128.820 595.700 133.820 596.820 ;
        RECT 135.540 595.700 137.180 596.820 ;
        RECT 138.900 595.700 143.900 596.820 ;
        RECT 145.620 595.700 150.620 596.820 ;
        RECT 152.340 595.700 157.340 596.820 ;
        RECT 159.060 595.700 160.700 596.820 ;
        RECT 162.420 595.700 167.420 596.820 ;
        RECT 169.140 595.700 174.140 596.820 ;
        RECT 175.860 595.700 177.500 596.820 ;
        RECT 179.220 595.700 184.220 596.820 ;
        RECT 185.940 595.700 190.940 596.820 ;
        RECT 192.660 595.700 197.660 596.820 ;
        RECT 199.380 595.700 201.020 596.820 ;
        RECT 202.740 595.700 207.740 596.820 ;
        RECT 209.460 595.700 214.460 596.820 ;
        RECT 216.180 595.700 217.820 596.820 ;
        RECT 219.540 595.700 224.540 596.820 ;
        RECT 226.260 595.700 231.260 596.820 ;
        RECT 232.980 595.700 237.980 596.820 ;
        RECT 239.700 595.700 241.340 596.820 ;
        RECT 243.060 595.700 248.060 596.820 ;
        RECT 249.780 595.700 254.780 596.820 ;
        RECT 256.500 595.700 261.500 596.820 ;
        RECT 263.220 595.700 264.860 596.820 ;
        RECT 266.580 595.700 271.580 596.820 ;
        RECT 273.300 595.700 278.300 596.820 ;
        RECT 280.020 595.700 281.660 596.820 ;
        RECT 283.380 595.700 288.380 596.820 ;
        RECT 290.100 595.700 295.100 596.820 ;
        RECT 296.820 595.700 301.820 596.820 ;
        RECT 303.540 595.700 305.180 596.820 ;
        RECT 306.900 595.700 311.900 596.820 ;
        RECT 313.620 595.700 318.620 596.820 ;
        RECT 320.340 595.700 325.340 596.820 ;
        RECT 327.060 595.700 328.700 596.820 ;
        RECT 330.420 595.700 335.420 596.820 ;
        RECT 337.140 595.700 342.140 596.820 ;
        RECT 343.860 595.700 345.500 596.820 ;
        RECT 347.220 595.700 352.220 596.820 ;
        RECT 353.940 595.700 358.940 596.820 ;
        RECT 360.660 595.700 365.660 596.820 ;
        RECT 367.380 595.700 369.020 596.820 ;
        RECT 370.740 595.700 375.740 596.820 ;
        RECT 377.460 595.700 382.460 596.820 ;
        RECT 384.180 595.700 389.180 596.820 ;
        RECT 390.900 595.700 392.540 596.820 ;
        RECT 394.260 595.700 399.260 596.820 ;
        RECT 400.980 595.700 405.980 596.820 ;
        RECT 407.700 595.700 409.340 596.820 ;
        RECT 411.060 595.700 416.060 596.820 ;
        RECT 417.780 595.700 422.780 596.820 ;
        RECT 424.500 595.700 429.500 596.820 ;
        RECT 431.220 595.700 432.860 596.820 ;
        RECT 434.580 595.700 439.580 596.820 ;
        RECT 441.300 595.700 446.300 596.820 ;
        RECT 448.020 595.700 453.020 596.820 ;
        RECT 454.740 595.700 456.380 596.820 ;
        RECT 458.100 595.700 463.100 596.820 ;
        RECT 464.820 595.700 469.820 596.820 ;
        RECT 471.540 595.700 473.180 596.820 ;
        RECT 474.900 595.700 479.900 596.820 ;
        RECT 481.620 595.700 486.620 596.820 ;
        RECT 488.340 595.700 493.340 596.820 ;
        RECT 495.060 595.700 496.700 596.820 ;
        RECT 498.420 595.700 503.420 596.820 ;
        RECT 505.140 595.700 510.140 596.820 ;
        RECT 511.860 595.700 513.500 596.820 ;
        RECT 515.220 595.700 520.220 596.820 ;
        RECT 521.940 595.700 526.940 596.820 ;
        RECT 528.660 595.700 533.660 596.820 ;
        RECT 535.380 595.700 537.020 596.820 ;
        RECT 538.740 595.700 543.740 596.820 ;
        RECT 545.460 595.700 550.460 596.820 ;
        RECT 552.180 595.700 557.180 596.820 ;
        RECT 558.900 595.700 560.540 596.820 ;
        RECT 562.260 595.700 567.260 596.820 ;
        RECT 568.980 595.700 573.980 596.820 ;
        RECT 575.700 595.700 577.340 596.820 ;
        RECT 579.060 595.700 584.060 596.820 ;
        RECT 585.780 595.700 590.780 596.820 ;
        RECT 592.500 595.700 594.580 596.820 ;
        RECT 0.700 4.300 594.580 595.700 ;
        RECT 1.140 3.500 2.780 4.300 ;
        RECT 4.500 3.500 9.500 4.300 ;
        RECT 11.220 3.500 16.220 4.300 ;
        RECT 17.940 3.500 19.580 4.300 ;
        RECT 21.300 3.500 26.300 4.300 ;
        RECT 28.020 3.500 33.020 4.300 ;
        RECT 34.740 3.500 39.740 4.300 ;
        RECT 41.460 3.500 43.100 4.300 ;
        RECT 44.820 3.500 49.820 4.300 ;
        RECT 51.540 3.500 56.540 4.300 ;
        RECT 58.260 3.500 59.900 4.300 ;
        RECT 61.620 3.500 66.620 4.300 ;
        RECT 68.340 3.500 73.340 4.300 ;
        RECT 75.060 3.500 80.060 4.300 ;
        RECT 81.780 3.500 83.420 4.300 ;
        RECT 85.140 3.500 90.140 4.300 ;
        RECT 91.860 3.500 96.860 4.300 ;
        RECT 98.580 3.500 103.580 4.300 ;
        RECT 105.300 3.500 106.940 4.300 ;
        RECT 108.660 3.500 113.660 4.300 ;
        RECT 115.380 3.500 120.380 4.300 ;
        RECT 122.100 3.500 123.740 4.300 ;
        RECT 125.460 3.500 130.460 4.300 ;
        RECT 132.180 3.500 137.180 4.300 ;
        RECT 138.900 3.500 143.900 4.300 ;
        RECT 145.620 3.500 147.260 4.300 ;
        RECT 148.980 3.500 153.980 4.300 ;
        RECT 155.700 3.500 160.700 4.300 ;
        RECT 162.420 3.500 167.420 4.300 ;
        RECT 169.140 3.500 170.780 4.300 ;
        RECT 172.500 3.500 177.500 4.300 ;
        RECT 179.220 3.500 184.220 4.300 ;
        RECT 185.940 3.500 187.580 4.300 ;
        RECT 189.300 3.500 194.300 4.300 ;
        RECT 196.020 3.500 201.020 4.300 ;
        RECT 202.740 3.500 207.740 4.300 ;
        RECT 209.460 3.500 211.100 4.300 ;
        RECT 212.820 3.500 217.820 4.300 ;
        RECT 219.540 3.500 224.540 4.300 ;
        RECT 226.260 3.500 231.260 4.300 ;
        RECT 232.980 3.500 234.620 4.300 ;
        RECT 236.340 3.500 241.340 4.300 ;
        RECT 243.060 3.500 248.060 4.300 ;
        RECT 249.780 3.500 251.420 4.300 ;
        RECT 253.140 3.500 258.140 4.300 ;
        RECT 259.860 3.500 264.860 4.300 ;
        RECT 266.580 3.500 271.580 4.300 ;
        RECT 273.300 3.500 274.940 4.300 ;
        RECT 276.660 3.500 281.660 4.300 ;
        RECT 283.380 3.500 288.380 4.300 ;
        RECT 290.100 3.500 291.740 4.300 ;
        RECT 293.460 3.500 298.460 4.300 ;
        RECT 300.180 3.500 305.180 4.300 ;
        RECT 306.900 3.500 311.900 4.300 ;
        RECT 313.620 3.500 315.260 4.300 ;
        RECT 316.980 3.500 321.980 4.300 ;
        RECT 323.700 3.500 328.700 4.300 ;
        RECT 330.420 3.500 335.420 4.300 ;
        RECT 337.140 3.500 338.780 4.300 ;
        RECT 340.500 3.500 345.500 4.300 ;
        RECT 347.220 3.500 352.220 4.300 ;
        RECT 353.940 3.500 355.580 4.300 ;
        RECT 357.300 3.500 362.300 4.300 ;
        RECT 364.020 3.500 369.020 4.300 ;
        RECT 370.740 3.500 375.740 4.300 ;
        RECT 377.460 3.500 379.100 4.300 ;
        RECT 380.820 3.500 385.820 4.300 ;
        RECT 387.540 3.500 392.540 4.300 ;
        RECT 394.260 3.500 399.260 4.300 ;
        RECT 400.980 3.500 402.620 4.300 ;
        RECT 404.340 3.500 409.340 4.300 ;
        RECT 411.060 3.500 416.060 4.300 ;
        RECT 417.780 3.500 419.420 4.300 ;
        RECT 421.140 3.500 426.140 4.300 ;
        RECT 427.860 3.500 432.860 4.300 ;
        RECT 434.580 3.500 439.580 4.300 ;
        RECT 441.300 3.500 442.940 4.300 ;
        RECT 444.660 3.500 449.660 4.300 ;
        RECT 451.380 3.500 456.380 4.300 ;
        RECT 458.100 3.500 463.100 4.300 ;
        RECT 464.820 3.500 466.460 4.300 ;
        RECT 468.180 3.500 473.180 4.300 ;
        RECT 474.900 3.500 479.900 4.300 ;
        RECT 481.620 3.500 483.260 4.300 ;
        RECT 484.980 3.500 489.980 4.300 ;
        RECT 491.700 3.500 496.700 4.300 ;
        RECT 498.420 3.500 503.420 4.300 ;
        RECT 505.140 3.500 506.780 4.300 ;
        RECT 508.500 3.500 513.500 4.300 ;
        RECT 515.220 3.500 520.220 4.300 ;
        RECT 521.940 3.500 526.940 4.300 ;
        RECT 528.660 3.500 530.300 4.300 ;
        RECT 532.020 3.500 537.020 4.300 ;
        RECT 538.740 3.500 543.740 4.300 ;
        RECT 545.460 3.500 547.100 4.300 ;
        RECT 548.820 3.500 553.820 4.300 ;
        RECT 555.540 3.500 560.540 4.300 ;
        RECT 562.260 3.500 567.260 4.300 ;
        RECT 568.980 3.500 570.620 4.300 ;
        RECT 572.340 3.500 577.340 4.300 ;
        RECT 579.060 3.500 584.060 4.300 ;
        RECT 585.780 3.500 587.420 4.300 ;
        RECT 589.140 3.500 594.140 4.300 ;
      LAYER Metal3 ;
        RECT 0.650 594.140 0.700 594.580 ;
        RECT 4.300 594.140 596.820 594.580 ;
        RECT 0.650 592.500 596.820 594.140 ;
        RECT 0.650 590.780 595.700 592.500 ;
        RECT 0.650 589.140 596.820 590.780 ;
        RECT 0.650 587.420 0.700 589.140 ;
        RECT 4.300 587.420 596.820 589.140 ;
        RECT 0.650 585.780 596.820 587.420 ;
        RECT 0.650 584.060 0.700 585.780 ;
        RECT 4.300 584.060 595.700 585.780 ;
        RECT 0.650 579.060 596.820 584.060 ;
        RECT 0.650 577.340 0.700 579.060 ;
        RECT 4.300 577.340 595.700 579.060 ;
        RECT 0.650 575.700 596.820 577.340 ;
        RECT 0.650 573.980 595.700 575.700 ;
        RECT 0.650 572.340 596.820 573.980 ;
        RECT 0.650 570.620 0.700 572.340 ;
        RECT 4.300 570.620 596.820 572.340 ;
        RECT 0.650 568.980 596.820 570.620 ;
        RECT 0.650 567.260 0.700 568.980 ;
        RECT 4.300 567.260 595.700 568.980 ;
        RECT 0.650 562.260 596.820 567.260 ;
        RECT 0.650 560.540 0.700 562.260 ;
        RECT 4.300 560.540 595.700 562.260 ;
        RECT 0.650 558.900 596.820 560.540 ;
        RECT 0.650 557.180 595.700 558.900 ;
        RECT 0.650 555.540 596.820 557.180 ;
        RECT 0.650 553.820 0.700 555.540 ;
        RECT 4.300 553.820 596.820 555.540 ;
        RECT 0.650 552.180 596.820 553.820 ;
        RECT 0.650 550.460 595.700 552.180 ;
        RECT 0.650 548.820 596.820 550.460 ;
        RECT 0.650 547.100 0.700 548.820 ;
        RECT 4.300 547.100 596.820 548.820 ;
        RECT 0.650 545.460 596.820 547.100 ;
        RECT 0.650 543.740 0.700 545.460 ;
        RECT 4.300 543.740 595.700 545.460 ;
        RECT 0.650 538.740 596.820 543.740 ;
        RECT 0.650 537.020 0.700 538.740 ;
        RECT 4.300 537.020 595.700 538.740 ;
        RECT 0.650 535.380 596.820 537.020 ;
        RECT 0.650 533.660 595.700 535.380 ;
        RECT 0.650 532.020 596.820 533.660 ;
        RECT 0.650 530.300 0.700 532.020 ;
        RECT 4.300 530.300 596.820 532.020 ;
        RECT 0.650 528.660 596.820 530.300 ;
        RECT 0.650 526.940 0.700 528.660 ;
        RECT 4.300 526.940 595.700 528.660 ;
        RECT 0.650 521.940 596.820 526.940 ;
        RECT 0.650 520.220 0.700 521.940 ;
        RECT 4.300 520.220 595.700 521.940 ;
        RECT 0.650 515.220 596.820 520.220 ;
        RECT 0.650 513.500 0.700 515.220 ;
        RECT 4.300 513.500 595.700 515.220 ;
        RECT 0.650 511.860 596.820 513.500 ;
        RECT 0.650 510.140 595.700 511.860 ;
        RECT 0.650 508.500 596.820 510.140 ;
        RECT 0.650 506.780 0.700 508.500 ;
        RECT 4.300 506.780 596.820 508.500 ;
        RECT 0.650 505.140 596.820 506.780 ;
        RECT 0.650 503.420 0.700 505.140 ;
        RECT 4.300 503.420 595.700 505.140 ;
        RECT 0.650 498.420 596.820 503.420 ;
        RECT 0.650 496.700 0.700 498.420 ;
        RECT 4.300 496.700 595.700 498.420 ;
        RECT 0.650 495.060 596.820 496.700 ;
        RECT 0.650 493.340 595.700 495.060 ;
        RECT 0.650 491.700 596.820 493.340 ;
        RECT 0.650 489.980 0.700 491.700 ;
        RECT 4.300 489.980 596.820 491.700 ;
        RECT 0.650 488.340 596.820 489.980 ;
        RECT 0.650 486.620 595.700 488.340 ;
        RECT 0.650 484.980 596.820 486.620 ;
        RECT 0.650 483.260 0.700 484.980 ;
        RECT 4.300 483.260 596.820 484.980 ;
        RECT 0.650 481.620 596.820 483.260 ;
        RECT 0.650 479.900 0.700 481.620 ;
        RECT 4.300 479.900 595.700 481.620 ;
        RECT 0.650 474.900 596.820 479.900 ;
        RECT 0.650 473.180 0.700 474.900 ;
        RECT 4.300 473.180 595.700 474.900 ;
        RECT 0.650 471.540 596.820 473.180 ;
        RECT 0.650 469.820 595.700 471.540 ;
        RECT 0.650 468.180 596.820 469.820 ;
        RECT 0.650 466.460 0.700 468.180 ;
        RECT 4.300 466.460 596.820 468.180 ;
        RECT 0.650 464.820 596.820 466.460 ;
        RECT 0.650 463.100 0.700 464.820 ;
        RECT 4.300 463.100 595.700 464.820 ;
        RECT 0.650 458.100 596.820 463.100 ;
        RECT 0.650 456.380 0.700 458.100 ;
        RECT 4.300 456.380 595.700 458.100 ;
        RECT 0.650 454.740 596.820 456.380 ;
        RECT 0.650 453.020 595.700 454.740 ;
        RECT 0.650 451.380 596.820 453.020 ;
        RECT 0.650 449.660 0.700 451.380 ;
        RECT 4.300 449.660 596.820 451.380 ;
        RECT 0.650 448.020 596.820 449.660 ;
        RECT 0.650 446.300 595.700 448.020 ;
        RECT 0.650 444.660 596.820 446.300 ;
        RECT 0.650 442.940 0.700 444.660 ;
        RECT 4.300 442.940 596.820 444.660 ;
        RECT 0.650 441.300 596.820 442.940 ;
        RECT 0.650 439.580 0.700 441.300 ;
        RECT 4.300 439.580 595.700 441.300 ;
        RECT 0.650 434.580 596.820 439.580 ;
        RECT 0.650 432.860 0.700 434.580 ;
        RECT 4.300 432.860 595.700 434.580 ;
        RECT 0.650 431.220 596.820 432.860 ;
        RECT 0.650 429.500 595.700 431.220 ;
        RECT 0.650 427.860 596.820 429.500 ;
        RECT 0.650 426.140 0.700 427.860 ;
        RECT 4.300 426.140 596.820 427.860 ;
        RECT 0.650 424.500 596.820 426.140 ;
        RECT 0.650 422.780 595.700 424.500 ;
        RECT 0.650 421.140 596.820 422.780 ;
        RECT 0.650 419.420 0.700 421.140 ;
        RECT 4.300 419.420 596.820 421.140 ;
        RECT 0.650 417.780 596.820 419.420 ;
        RECT 0.650 416.060 0.700 417.780 ;
        RECT 4.300 416.060 595.700 417.780 ;
        RECT 0.650 411.060 596.820 416.060 ;
        RECT 0.650 409.340 0.700 411.060 ;
        RECT 4.300 409.340 595.700 411.060 ;
        RECT 0.650 407.700 596.820 409.340 ;
        RECT 0.650 405.980 595.700 407.700 ;
        RECT 0.650 404.340 596.820 405.980 ;
        RECT 0.650 402.620 0.700 404.340 ;
        RECT 4.300 402.620 596.820 404.340 ;
        RECT 0.650 400.980 596.820 402.620 ;
        RECT 0.650 399.260 0.700 400.980 ;
        RECT 4.300 399.260 595.700 400.980 ;
        RECT 0.650 394.260 596.820 399.260 ;
        RECT 0.650 392.540 0.700 394.260 ;
        RECT 4.300 392.540 595.700 394.260 ;
        RECT 0.650 390.900 596.820 392.540 ;
        RECT 0.650 389.180 595.700 390.900 ;
        RECT 0.650 387.540 596.820 389.180 ;
        RECT 0.650 385.820 0.700 387.540 ;
        RECT 4.300 385.820 596.820 387.540 ;
        RECT 0.650 384.180 596.820 385.820 ;
        RECT 0.650 382.460 595.700 384.180 ;
        RECT 0.650 380.820 596.820 382.460 ;
        RECT 0.650 379.100 0.700 380.820 ;
        RECT 4.300 379.100 596.820 380.820 ;
        RECT 0.650 377.460 596.820 379.100 ;
        RECT 0.650 375.740 0.700 377.460 ;
        RECT 4.300 375.740 595.700 377.460 ;
        RECT 0.650 370.740 596.820 375.740 ;
        RECT 0.650 369.020 0.700 370.740 ;
        RECT 4.300 369.020 595.700 370.740 ;
        RECT 0.650 367.380 596.820 369.020 ;
        RECT 0.650 365.660 595.700 367.380 ;
        RECT 0.650 364.020 596.820 365.660 ;
        RECT 0.650 362.300 0.700 364.020 ;
        RECT 4.300 362.300 596.820 364.020 ;
        RECT 0.650 360.660 596.820 362.300 ;
        RECT 0.650 358.940 595.700 360.660 ;
        RECT 0.650 357.300 596.820 358.940 ;
        RECT 0.650 355.580 0.700 357.300 ;
        RECT 4.300 355.580 596.820 357.300 ;
        RECT 0.650 353.940 596.820 355.580 ;
        RECT 0.650 352.220 0.700 353.940 ;
        RECT 4.300 352.220 595.700 353.940 ;
        RECT 0.650 347.220 596.820 352.220 ;
        RECT 0.650 345.500 0.700 347.220 ;
        RECT 4.300 345.500 595.700 347.220 ;
        RECT 0.650 343.860 596.820 345.500 ;
        RECT 0.650 342.140 595.700 343.860 ;
        RECT 0.650 340.500 596.820 342.140 ;
        RECT 0.650 338.780 0.700 340.500 ;
        RECT 4.300 338.780 596.820 340.500 ;
        RECT 0.650 337.140 596.820 338.780 ;
        RECT 0.650 335.420 0.700 337.140 ;
        RECT 4.300 335.420 595.700 337.140 ;
        RECT 0.650 330.420 596.820 335.420 ;
        RECT 0.650 328.700 0.700 330.420 ;
        RECT 4.300 328.700 595.700 330.420 ;
        RECT 0.650 327.060 596.820 328.700 ;
        RECT 0.650 325.340 595.700 327.060 ;
        RECT 0.650 323.700 596.820 325.340 ;
        RECT 0.650 321.980 0.700 323.700 ;
        RECT 4.300 321.980 596.820 323.700 ;
        RECT 0.650 320.340 596.820 321.980 ;
        RECT 0.650 318.620 595.700 320.340 ;
        RECT 0.650 316.980 596.820 318.620 ;
        RECT 0.650 315.260 0.700 316.980 ;
        RECT 4.300 315.260 596.820 316.980 ;
        RECT 0.650 313.620 596.820 315.260 ;
        RECT 0.650 311.900 0.700 313.620 ;
        RECT 4.300 311.900 595.700 313.620 ;
        RECT 0.650 306.900 596.820 311.900 ;
        RECT 0.650 305.180 0.700 306.900 ;
        RECT 4.300 305.180 595.700 306.900 ;
        RECT 0.650 303.540 596.820 305.180 ;
        RECT 0.650 301.820 595.700 303.540 ;
        RECT 0.650 300.180 596.820 301.820 ;
        RECT 0.650 298.460 0.700 300.180 ;
        RECT 4.300 298.460 596.820 300.180 ;
        RECT 0.650 296.820 596.820 298.460 ;
        RECT 0.650 295.100 595.700 296.820 ;
        RECT 0.650 293.460 596.820 295.100 ;
        RECT 0.650 291.740 0.700 293.460 ;
        RECT 4.300 291.740 596.820 293.460 ;
        RECT 0.650 290.100 596.820 291.740 ;
        RECT 0.650 288.380 0.700 290.100 ;
        RECT 4.300 288.380 595.700 290.100 ;
        RECT 0.650 283.380 596.820 288.380 ;
        RECT 0.650 281.660 0.700 283.380 ;
        RECT 4.300 281.660 595.700 283.380 ;
        RECT 0.650 280.020 596.820 281.660 ;
        RECT 0.650 278.300 595.700 280.020 ;
        RECT 0.650 276.660 596.820 278.300 ;
        RECT 0.650 274.940 0.700 276.660 ;
        RECT 4.300 274.940 596.820 276.660 ;
        RECT 0.650 273.300 596.820 274.940 ;
        RECT 0.650 271.580 0.700 273.300 ;
        RECT 4.300 271.580 595.700 273.300 ;
        RECT 0.650 266.580 596.820 271.580 ;
        RECT 0.650 264.860 0.700 266.580 ;
        RECT 4.300 264.860 595.700 266.580 ;
        RECT 0.650 263.220 596.820 264.860 ;
        RECT 0.650 261.500 595.700 263.220 ;
        RECT 0.650 259.860 596.820 261.500 ;
        RECT 0.650 258.140 0.700 259.860 ;
        RECT 4.300 258.140 596.820 259.860 ;
        RECT 0.650 256.500 596.820 258.140 ;
        RECT 0.650 254.780 595.700 256.500 ;
        RECT 0.650 253.140 596.820 254.780 ;
        RECT 0.650 251.420 0.700 253.140 ;
        RECT 4.300 251.420 596.820 253.140 ;
        RECT 0.650 249.780 596.820 251.420 ;
        RECT 0.650 248.060 0.700 249.780 ;
        RECT 4.300 248.060 595.700 249.780 ;
        RECT 0.650 243.060 596.820 248.060 ;
        RECT 0.650 241.340 0.700 243.060 ;
        RECT 4.300 241.340 595.700 243.060 ;
        RECT 0.650 239.700 596.820 241.340 ;
        RECT 0.650 237.980 595.700 239.700 ;
        RECT 0.650 236.340 596.820 237.980 ;
        RECT 0.650 234.620 0.700 236.340 ;
        RECT 4.300 234.620 596.820 236.340 ;
        RECT 0.650 232.980 596.820 234.620 ;
        RECT 0.650 231.260 0.700 232.980 ;
        RECT 4.300 231.260 595.700 232.980 ;
        RECT 0.650 226.260 596.820 231.260 ;
        RECT 0.650 224.540 0.700 226.260 ;
        RECT 4.300 224.540 595.700 226.260 ;
        RECT 0.650 219.540 596.820 224.540 ;
        RECT 0.650 217.820 0.700 219.540 ;
        RECT 4.300 217.820 595.700 219.540 ;
        RECT 0.650 216.180 596.820 217.820 ;
        RECT 0.650 214.460 595.700 216.180 ;
        RECT 0.650 212.820 596.820 214.460 ;
        RECT 0.650 211.100 0.700 212.820 ;
        RECT 4.300 211.100 596.820 212.820 ;
        RECT 0.650 209.460 596.820 211.100 ;
        RECT 0.650 207.740 0.700 209.460 ;
        RECT 4.300 207.740 595.700 209.460 ;
        RECT 0.650 202.740 596.820 207.740 ;
        RECT 0.650 201.020 0.700 202.740 ;
        RECT 4.300 201.020 595.700 202.740 ;
        RECT 0.650 199.380 596.820 201.020 ;
        RECT 0.650 197.660 595.700 199.380 ;
        RECT 0.650 196.020 596.820 197.660 ;
        RECT 0.650 194.300 0.700 196.020 ;
        RECT 4.300 194.300 596.820 196.020 ;
        RECT 0.650 192.660 596.820 194.300 ;
        RECT 0.650 190.940 595.700 192.660 ;
        RECT 0.650 189.300 596.820 190.940 ;
        RECT 0.650 187.580 0.700 189.300 ;
        RECT 4.300 187.580 596.820 189.300 ;
        RECT 0.650 185.940 596.820 187.580 ;
        RECT 0.650 184.220 0.700 185.940 ;
        RECT 4.300 184.220 595.700 185.940 ;
        RECT 0.650 179.220 596.820 184.220 ;
        RECT 0.650 177.500 0.700 179.220 ;
        RECT 4.300 177.500 595.700 179.220 ;
        RECT 0.650 175.860 596.820 177.500 ;
        RECT 0.650 174.140 595.700 175.860 ;
        RECT 0.650 172.500 596.820 174.140 ;
        RECT 0.650 170.780 0.700 172.500 ;
        RECT 4.300 170.780 596.820 172.500 ;
        RECT 0.650 169.140 596.820 170.780 ;
        RECT 0.650 167.420 0.700 169.140 ;
        RECT 4.300 167.420 595.700 169.140 ;
        RECT 0.650 162.420 596.820 167.420 ;
        RECT 0.650 160.700 0.700 162.420 ;
        RECT 4.300 160.700 595.700 162.420 ;
        RECT 0.650 159.060 596.820 160.700 ;
        RECT 0.650 157.340 595.700 159.060 ;
        RECT 0.650 155.700 596.820 157.340 ;
        RECT 0.650 153.980 0.700 155.700 ;
        RECT 4.300 153.980 596.820 155.700 ;
        RECT 0.650 152.340 596.820 153.980 ;
        RECT 0.650 150.620 595.700 152.340 ;
        RECT 0.650 148.980 596.820 150.620 ;
        RECT 0.650 147.260 0.700 148.980 ;
        RECT 4.300 147.260 596.820 148.980 ;
        RECT 0.650 145.620 596.820 147.260 ;
        RECT 0.650 143.900 0.700 145.620 ;
        RECT 4.300 143.900 595.700 145.620 ;
        RECT 0.650 138.900 596.820 143.900 ;
        RECT 0.650 137.180 0.700 138.900 ;
        RECT 4.300 137.180 595.700 138.900 ;
        RECT 0.650 135.540 596.820 137.180 ;
        RECT 0.650 133.820 595.700 135.540 ;
        RECT 0.650 132.180 596.820 133.820 ;
        RECT 0.650 130.460 0.700 132.180 ;
        RECT 4.300 130.460 596.820 132.180 ;
        RECT 0.650 128.820 596.820 130.460 ;
        RECT 0.650 127.100 595.700 128.820 ;
        RECT 0.650 125.460 596.820 127.100 ;
        RECT 0.650 123.740 0.700 125.460 ;
        RECT 4.300 123.740 596.820 125.460 ;
        RECT 0.650 122.100 596.820 123.740 ;
        RECT 0.650 120.380 0.700 122.100 ;
        RECT 4.300 120.380 595.700 122.100 ;
        RECT 0.650 115.380 596.820 120.380 ;
        RECT 0.650 113.660 0.700 115.380 ;
        RECT 4.300 113.660 595.700 115.380 ;
        RECT 0.650 112.020 596.820 113.660 ;
        RECT 0.650 110.300 595.700 112.020 ;
        RECT 0.650 108.660 596.820 110.300 ;
        RECT 0.650 106.940 0.700 108.660 ;
        RECT 4.300 106.940 596.820 108.660 ;
        RECT 0.650 105.300 596.820 106.940 ;
        RECT 0.650 103.580 0.700 105.300 ;
        RECT 4.300 103.580 595.700 105.300 ;
        RECT 0.650 98.580 596.820 103.580 ;
        RECT 0.650 96.860 0.700 98.580 ;
        RECT 4.300 96.860 595.700 98.580 ;
        RECT 0.650 95.220 596.820 96.860 ;
        RECT 0.650 93.500 595.700 95.220 ;
        RECT 0.650 91.860 596.820 93.500 ;
        RECT 0.650 90.140 0.700 91.860 ;
        RECT 4.300 90.140 596.820 91.860 ;
        RECT 0.650 88.500 596.820 90.140 ;
        RECT 0.650 86.780 595.700 88.500 ;
        RECT 0.650 85.140 596.820 86.780 ;
        RECT 0.650 83.420 0.700 85.140 ;
        RECT 4.300 83.420 596.820 85.140 ;
        RECT 0.650 81.780 596.820 83.420 ;
        RECT 0.650 80.060 0.700 81.780 ;
        RECT 4.300 80.060 595.700 81.780 ;
        RECT 0.650 75.060 596.820 80.060 ;
        RECT 0.650 73.340 0.700 75.060 ;
        RECT 4.300 73.340 595.700 75.060 ;
        RECT 0.650 71.700 596.820 73.340 ;
        RECT 0.650 69.980 595.700 71.700 ;
        RECT 0.650 68.340 596.820 69.980 ;
        RECT 0.650 66.620 0.700 68.340 ;
        RECT 4.300 66.620 596.820 68.340 ;
        RECT 0.650 64.980 596.820 66.620 ;
        RECT 0.650 63.260 595.700 64.980 ;
        RECT 0.650 61.620 596.820 63.260 ;
        RECT 0.650 59.900 0.700 61.620 ;
        RECT 4.300 59.900 596.820 61.620 ;
        RECT 0.650 58.260 596.820 59.900 ;
        RECT 0.650 56.540 0.700 58.260 ;
        RECT 4.300 56.540 595.700 58.260 ;
        RECT 0.650 51.540 596.820 56.540 ;
        RECT 0.650 49.820 0.700 51.540 ;
        RECT 4.300 49.820 595.700 51.540 ;
        RECT 0.650 48.180 596.820 49.820 ;
        RECT 0.650 46.460 595.700 48.180 ;
        RECT 0.650 44.820 596.820 46.460 ;
        RECT 0.650 43.100 0.700 44.820 ;
        RECT 4.300 43.100 596.820 44.820 ;
        RECT 0.650 41.460 596.820 43.100 ;
        RECT 0.650 39.740 0.700 41.460 ;
        RECT 4.300 39.740 595.700 41.460 ;
        RECT 0.650 34.740 596.820 39.740 ;
        RECT 0.650 33.020 0.700 34.740 ;
        RECT 4.300 33.020 595.700 34.740 ;
        RECT 0.650 31.380 596.820 33.020 ;
        RECT 0.650 29.660 595.700 31.380 ;
        RECT 0.650 28.020 596.820 29.660 ;
        RECT 0.650 26.300 0.700 28.020 ;
        RECT 4.300 26.300 596.820 28.020 ;
        RECT 0.650 24.660 596.820 26.300 ;
        RECT 0.650 22.940 595.700 24.660 ;
        RECT 0.650 21.300 596.820 22.940 ;
        RECT 0.650 19.580 0.700 21.300 ;
        RECT 4.300 19.580 596.820 21.300 ;
        RECT 0.650 17.940 596.820 19.580 ;
        RECT 0.650 16.220 0.700 17.940 ;
        RECT 4.300 16.220 595.700 17.940 ;
        RECT 0.650 11.220 596.820 16.220 ;
        RECT 0.650 9.500 0.700 11.220 ;
        RECT 4.300 9.500 595.700 11.220 ;
        RECT 0.650 7.860 596.820 9.500 ;
        RECT 0.650 7.420 595.700 7.860 ;
      LAYER Metal4 ;
        RECT 238.700 218.490 252.340 316.870 ;
        RECT 254.540 218.490 329.140 316.870 ;
        RECT 331.340 218.490 366.660 316.870 ;
  END
END user_proj_example
END LIBRARY

