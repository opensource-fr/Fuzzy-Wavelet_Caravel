magic
tech gf180mcuC
magscale 1 5
timestamp 1670287222
<< obsm1 >>
rect 672 855 59304 58561
<< metal2 >>
rect -28 59600 84 59900
rect 644 59600 756 59900
rect 980 59600 1092 59900
rect 1652 59600 1764 59900
rect 2324 59600 2436 59900
rect 2996 59600 3108 59900
rect 3332 59600 3444 59900
rect 4004 59600 4116 59900
rect 4676 59600 4788 59900
rect 5012 59600 5124 59900
rect 5684 59600 5796 59900
rect 6356 59600 6468 59900
rect 7028 59600 7140 59900
rect 7364 59600 7476 59900
rect 8036 59600 8148 59900
rect 8708 59600 8820 59900
rect 9380 59600 9492 59900
rect 9716 59600 9828 59900
rect 10388 59600 10500 59900
rect 11060 59600 11172 59900
rect 11396 59600 11508 59900
rect 12068 59600 12180 59900
rect 12740 59600 12852 59900
rect 13412 59600 13524 59900
rect 13748 59600 13860 59900
rect 14420 59600 14532 59900
rect 15092 59600 15204 59900
rect 15764 59600 15876 59900
rect 16100 59600 16212 59900
rect 16772 59600 16884 59900
rect 17444 59600 17556 59900
rect 17780 59600 17892 59900
rect 18452 59600 18564 59900
rect 19124 59600 19236 59900
rect 19796 59600 19908 59900
rect 20132 59600 20244 59900
rect 20804 59600 20916 59900
rect 21476 59600 21588 59900
rect 21812 59600 21924 59900
rect 22484 59600 22596 59900
rect 23156 59600 23268 59900
rect 23828 59600 23940 59900
rect 24164 59600 24276 59900
rect 24836 59600 24948 59900
rect 25508 59600 25620 59900
rect 26180 59600 26292 59900
rect 26516 59600 26628 59900
rect 27188 59600 27300 59900
rect 27860 59600 27972 59900
rect 28196 59600 28308 59900
rect 28868 59600 28980 59900
rect 29540 59600 29652 59900
rect 30212 59600 30324 59900
rect 30548 59600 30660 59900
rect 31220 59600 31332 59900
rect 31892 59600 32004 59900
rect 32564 59600 32676 59900
rect 32900 59600 33012 59900
rect 33572 59600 33684 59900
rect 34244 59600 34356 59900
rect 34580 59600 34692 59900
rect 35252 59600 35364 59900
rect 35924 59600 36036 59900
rect 36596 59600 36708 59900
rect 36932 59600 37044 59900
rect 37604 59600 37716 59900
rect 38276 59600 38388 59900
rect 38948 59600 39060 59900
rect 39284 59600 39396 59900
rect 39956 59600 40068 59900
rect 40628 59600 40740 59900
rect 40964 59600 41076 59900
rect 41636 59600 41748 59900
rect 42308 59600 42420 59900
rect 42980 59600 43092 59900
rect 43316 59600 43428 59900
rect 43988 59600 44100 59900
rect 44660 59600 44772 59900
rect 45332 59600 45444 59900
rect 45668 59600 45780 59900
rect 46340 59600 46452 59900
rect 47012 59600 47124 59900
rect 47348 59600 47460 59900
rect 48020 59600 48132 59900
rect 48692 59600 48804 59900
rect 49364 59600 49476 59900
rect 49700 59600 49812 59900
rect 50372 59600 50484 59900
rect 51044 59600 51156 59900
rect 51380 59600 51492 59900
rect 52052 59600 52164 59900
rect 52724 59600 52836 59900
rect 53396 59600 53508 59900
rect 53732 59600 53844 59900
rect 54404 59600 54516 59900
rect 55076 59600 55188 59900
rect 55748 59600 55860 59900
rect 56084 59600 56196 59900
rect 56756 59600 56868 59900
rect 57428 59600 57540 59900
rect 57764 59600 57876 59900
rect 58436 59600 58548 59900
rect 59108 59600 59220 59900
rect 59780 59600 59892 59900
rect -28 100 84 400
rect 308 100 420 400
rect 980 100 1092 400
rect 1652 100 1764 400
rect 1988 100 2100 400
rect 2660 100 2772 400
rect 3332 100 3444 400
rect 4004 100 4116 400
rect 4340 100 4452 400
rect 5012 100 5124 400
rect 5684 100 5796 400
rect 6020 100 6132 400
rect 6692 100 6804 400
rect 7364 100 7476 400
rect 8036 100 8148 400
rect 8372 100 8484 400
rect 9044 100 9156 400
rect 9716 100 9828 400
rect 10388 100 10500 400
rect 10724 100 10836 400
rect 11396 100 11508 400
rect 12068 100 12180 400
rect 12404 100 12516 400
rect 13076 100 13188 400
rect 13748 100 13860 400
rect 14420 100 14532 400
rect 14756 100 14868 400
rect 15428 100 15540 400
rect 16100 100 16212 400
rect 16772 100 16884 400
rect 17108 100 17220 400
rect 17780 100 17892 400
rect 18452 100 18564 400
rect 18788 100 18900 400
rect 19460 100 19572 400
rect 20132 100 20244 400
rect 20804 100 20916 400
rect 21140 100 21252 400
rect 21812 100 21924 400
rect 22484 100 22596 400
rect 23156 100 23268 400
rect 23492 100 23604 400
rect 24164 100 24276 400
rect 24836 100 24948 400
rect 25172 100 25284 400
rect 25844 100 25956 400
rect 26516 100 26628 400
rect 27188 100 27300 400
rect 27524 100 27636 400
rect 28196 100 28308 400
rect 28868 100 28980 400
rect 29204 100 29316 400
rect 29876 100 29988 400
rect 30548 100 30660 400
rect 31220 100 31332 400
rect 31556 100 31668 400
rect 32228 100 32340 400
rect 32900 100 33012 400
rect 33572 100 33684 400
rect 33908 100 34020 400
rect 34580 100 34692 400
rect 35252 100 35364 400
rect 35588 100 35700 400
rect 36260 100 36372 400
rect 36932 100 37044 400
rect 37604 100 37716 400
rect 37940 100 38052 400
rect 38612 100 38724 400
rect 39284 100 39396 400
rect 39956 100 40068 400
rect 40292 100 40404 400
rect 40964 100 41076 400
rect 41636 100 41748 400
rect 41972 100 42084 400
rect 42644 100 42756 400
rect 43316 100 43428 400
rect 43988 100 44100 400
rect 44324 100 44436 400
rect 44996 100 45108 400
rect 45668 100 45780 400
rect 46340 100 46452 400
rect 46676 100 46788 400
rect 47348 100 47460 400
rect 48020 100 48132 400
rect 48356 100 48468 400
rect 49028 100 49140 400
rect 49700 100 49812 400
rect 50372 100 50484 400
rect 50708 100 50820 400
rect 51380 100 51492 400
rect 52052 100 52164 400
rect 52724 100 52836 400
rect 53060 100 53172 400
rect 53732 100 53844 400
rect 54404 100 54516 400
rect 54740 100 54852 400
rect 55412 100 55524 400
rect 56084 100 56196 400
rect 56756 100 56868 400
rect 57092 100 57204 400
rect 57764 100 57876 400
rect 58436 100 58548 400
rect 58772 100 58884 400
rect 59444 100 59556 400
<< obsm2 >>
rect 114 59570 614 59682
rect 786 59570 950 59682
rect 1122 59570 1622 59682
rect 1794 59570 2294 59682
rect 2466 59570 2966 59682
rect 3138 59570 3302 59682
rect 3474 59570 3974 59682
rect 4146 59570 4646 59682
rect 4818 59570 4982 59682
rect 5154 59570 5654 59682
rect 5826 59570 6326 59682
rect 6498 59570 6998 59682
rect 7170 59570 7334 59682
rect 7506 59570 8006 59682
rect 8178 59570 8678 59682
rect 8850 59570 9350 59682
rect 9522 59570 9686 59682
rect 9858 59570 10358 59682
rect 10530 59570 11030 59682
rect 11202 59570 11366 59682
rect 11538 59570 12038 59682
rect 12210 59570 12710 59682
rect 12882 59570 13382 59682
rect 13554 59570 13718 59682
rect 13890 59570 14390 59682
rect 14562 59570 15062 59682
rect 15234 59570 15734 59682
rect 15906 59570 16070 59682
rect 16242 59570 16742 59682
rect 16914 59570 17414 59682
rect 17586 59570 17750 59682
rect 17922 59570 18422 59682
rect 18594 59570 19094 59682
rect 19266 59570 19766 59682
rect 19938 59570 20102 59682
rect 20274 59570 20774 59682
rect 20946 59570 21446 59682
rect 21618 59570 21782 59682
rect 21954 59570 22454 59682
rect 22626 59570 23126 59682
rect 23298 59570 23798 59682
rect 23970 59570 24134 59682
rect 24306 59570 24806 59682
rect 24978 59570 25478 59682
rect 25650 59570 26150 59682
rect 26322 59570 26486 59682
rect 26658 59570 27158 59682
rect 27330 59570 27830 59682
rect 28002 59570 28166 59682
rect 28338 59570 28838 59682
rect 29010 59570 29510 59682
rect 29682 59570 30182 59682
rect 30354 59570 30518 59682
rect 30690 59570 31190 59682
rect 31362 59570 31862 59682
rect 32034 59570 32534 59682
rect 32706 59570 32870 59682
rect 33042 59570 33542 59682
rect 33714 59570 34214 59682
rect 34386 59570 34550 59682
rect 34722 59570 35222 59682
rect 35394 59570 35894 59682
rect 36066 59570 36566 59682
rect 36738 59570 36902 59682
rect 37074 59570 37574 59682
rect 37746 59570 38246 59682
rect 38418 59570 38918 59682
rect 39090 59570 39254 59682
rect 39426 59570 39926 59682
rect 40098 59570 40598 59682
rect 40770 59570 40934 59682
rect 41106 59570 41606 59682
rect 41778 59570 42278 59682
rect 42450 59570 42950 59682
rect 43122 59570 43286 59682
rect 43458 59570 43958 59682
rect 44130 59570 44630 59682
rect 44802 59570 45302 59682
rect 45474 59570 45638 59682
rect 45810 59570 46310 59682
rect 46482 59570 46982 59682
rect 47154 59570 47318 59682
rect 47490 59570 47990 59682
rect 48162 59570 48662 59682
rect 48834 59570 49334 59682
rect 49506 59570 49670 59682
rect 49842 59570 50342 59682
rect 50514 59570 51014 59682
rect 51186 59570 51350 59682
rect 51522 59570 52022 59682
rect 52194 59570 52694 59682
rect 52866 59570 53366 59682
rect 53538 59570 53702 59682
rect 53874 59570 54374 59682
rect 54546 59570 55046 59682
rect 55218 59570 55718 59682
rect 55890 59570 56054 59682
rect 56226 59570 56726 59682
rect 56898 59570 57398 59682
rect 57570 59570 57734 59682
rect 57906 59570 58406 59682
rect 58578 59570 59078 59682
rect 59250 59570 59458 59682
rect 70 430 59458 59570
rect 114 350 278 430
rect 450 350 950 430
rect 1122 350 1622 430
rect 1794 350 1958 430
rect 2130 350 2630 430
rect 2802 350 3302 430
rect 3474 350 3974 430
rect 4146 350 4310 430
rect 4482 350 4982 430
rect 5154 350 5654 430
rect 5826 350 5990 430
rect 6162 350 6662 430
rect 6834 350 7334 430
rect 7506 350 8006 430
rect 8178 350 8342 430
rect 8514 350 9014 430
rect 9186 350 9686 430
rect 9858 350 10358 430
rect 10530 350 10694 430
rect 10866 350 11366 430
rect 11538 350 12038 430
rect 12210 350 12374 430
rect 12546 350 13046 430
rect 13218 350 13718 430
rect 13890 350 14390 430
rect 14562 350 14726 430
rect 14898 350 15398 430
rect 15570 350 16070 430
rect 16242 350 16742 430
rect 16914 350 17078 430
rect 17250 350 17750 430
rect 17922 350 18422 430
rect 18594 350 18758 430
rect 18930 350 19430 430
rect 19602 350 20102 430
rect 20274 350 20774 430
rect 20946 350 21110 430
rect 21282 350 21782 430
rect 21954 350 22454 430
rect 22626 350 23126 430
rect 23298 350 23462 430
rect 23634 350 24134 430
rect 24306 350 24806 430
rect 24978 350 25142 430
rect 25314 350 25814 430
rect 25986 350 26486 430
rect 26658 350 27158 430
rect 27330 350 27494 430
rect 27666 350 28166 430
rect 28338 350 28838 430
rect 29010 350 29174 430
rect 29346 350 29846 430
rect 30018 350 30518 430
rect 30690 350 31190 430
rect 31362 350 31526 430
rect 31698 350 32198 430
rect 32370 350 32870 430
rect 33042 350 33542 430
rect 33714 350 33878 430
rect 34050 350 34550 430
rect 34722 350 35222 430
rect 35394 350 35558 430
rect 35730 350 36230 430
rect 36402 350 36902 430
rect 37074 350 37574 430
rect 37746 350 37910 430
rect 38082 350 38582 430
rect 38754 350 39254 430
rect 39426 350 39926 430
rect 40098 350 40262 430
rect 40434 350 40934 430
rect 41106 350 41606 430
rect 41778 350 41942 430
rect 42114 350 42614 430
rect 42786 350 43286 430
rect 43458 350 43958 430
rect 44130 350 44294 430
rect 44466 350 44966 430
rect 45138 350 45638 430
rect 45810 350 46310 430
rect 46482 350 46646 430
rect 46818 350 47318 430
rect 47490 350 47990 430
rect 48162 350 48326 430
rect 48498 350 48998 430
rect 49170 350 49670 430
rect 49842 350 50342 430
rect 50514 350 50678 430
rect 50850 350 51350 430
rect 51522 350 52022 430
rect 52194 350 52694 430
rect 52866 350 53030 430
rect 53202 350 53702 430
rect 53874 350 54374 430
rect 54546 350 54710 430
rect 54882 350 55382 430
rect 55554 350 56054 430
rect 56226 350 56726 430
rect 56898 350 57062 430
rect 57234 350 57734 430
rect 57906 350 58406 430
rect 58578 350 58742 430
rect 58914 350 59414 430
<< metal3 >>
rect 59600 59780 59900 59892
rect 100 59444 400 59556
rect 59600 59108 59900 59220
rect 100 58772 400 58884
rect 100 58436 400 58548
rect 59600 58436 59900 58548
rect 100 57764 400 57876
rect 59600 57764 59900 57876
rect 59600 57428 59900 57540
rect 100 57092 400 57204
rect 100 56756 400 56868
rect 59600 56756 59900 56868
rect 100 56084 400 56196
rect 59600 56084 59900 56196
rect 59600 55748 59900 55860
rect 100 55412 400 55524
rect 59600 55076 59900 55188
rect 100 54740 400 54852
rect 100 54404 400 54516
rect 59600 54404 59900 54516
rect 100 53732 400 53844
rect 59600 53732 59900 53844
rect 59600 53396 59900 53508
rect 100 53060 400 53172
rect 100 52724 400 52836
rect 59600 52724 59900 52836
rect 100 52052 400 52164
rect 59600 52052 59900 52164
rect 100 51380 400 51492
rect 59600 51380 59900 51492
rect 59600 51044 59900 51156
rect 100 50708 400 50820
rect 100 50372 400 50484
rect 59600 50372 59900 50484
rect 100 49700 400 49812
rect 59600 49700 59900 49812
rect 59600 49364 59900 49476
rect 100 49028 400 49140
rect 59600 48692 59900 48804
rect 100 48356 400 48468
rect 100 48020 400 48132
rect 59600 48020 59900 48132
rect 100 47348 400 47460
rect 59600 47348 59900 47460
rect 59600 47012 59900 47124
rect 100 46676 400 46788
rect 100 46340 400 46452
rect 59600 46340 59900 46452
rect 100 45668 400 45780
rect 59600 45668 59900 45780
rect 59600 45332 59900 45444
rect 100 44996 400 45108
rect 59600 44660 59900 44772
rect 100 44324 400 44436
rect 100 43988 400 44100
rect 59600 43988 59900 44100
rect 100 43316 400 43428
rect 59600 43316 59900 43428
rect 59600 42980 59900 43092
rect 100 42644 400 42756
rect 59600 42308 59900 42420
rect 100 41972 400 42084
rect 100 41636 400 41748
rect 59600 41636 59900 41748
rect 100 40964 400 41076
rect 59600 40964 59900 41076
rect 59600 40628 59900 40740
rect 100 40292 400 40404
rect 100 39956 400 40068
rect 59600 39956 59900 40068
rect 100 39284 400 39396
rect 59600 39284 59900 39396
rect 59600 38948 59900 39060
rect 100 38612 400 38724
rect 59600 38276 59900 38388
rect 100 37940 400 38052
rect 100 37604 400 37716
rect 59600 37604 59900 37716
rect 100 36932 400 37044
rect 59600 36932 59900 37044
rect 59600 36596 59900 36708
rect 100 36260 400 36372
rect 59600 35924 59900 36036
rect 100 35588 400 35700
rect 100 35252 400 35364
rect 59600 35252 59900 35364
rect 100 34580 400 34692
rect 59600 34580 59900 34692
rect 59600 34244 59900 34356
rect 100 33908 400 34020
rect 100 33572 400 33684
rect 59600 33572 59900 33684
rect 100 32900 400 33012
rect 59600 32900 59900 33012
rect 59600 32564 59900 32676
rect 100 32228 400 32340
rect 59600 31892 59900 32004
rect 100 31556 400 31668
rect 100 31220 400 31332
rect 59600 31220 59900 31332
rect 100 30548 400 30660
rect 59600 30548 59900 30660
rect 59600 30212 59900 30324
rect 100 29876 400 29988
rect 59600 29540 59900 29652
rect 100 29204 400 29316
rect 100 28868 400 28980
rect 59600 28868 59900 28980
rect 100 28196 400 28308
rect 59600 28196 59900 28308
rect 59600 27860 59900 27972
rect 100 27524 400 27636
rect 100 27188 400 27300
rect 59600 27188 59900 27300
rect 100 26516 400 26628
rect 59600 26516 59900 26628
rect 59600 26180 59900 26292
rect 100 25844 400 25956
rect 59600 25508 59900 25620
rect 100 25172 400 25284
rect 100 24836 400 24948
rect 59600 24836 59900 24948
rect 100 24164 400 24276
rect 59600 24164 59900 24276
rect 59600 23828 59900 23940
rect 100 23492 400 23604
rect 100 23156 400 23268
rect 59600 23156 59900 23268
rect 100 22484 400 22596
rect 59600 22484 59900 22596
rect 100 21812 400 21924
rect 59600 21812 59900 21924
rect 59600 21476 59900 21588
rect 100 21140 400 21252
rect 100 20804 400 20916
rect 59600 20804 59900 20916
rect 100 20132 400 20244
rect 59600 20132 59900 20244
rect 59600 19796 59900 19908
rect 100 19460 400 19572
rect 59600 19124 59900 19236
rect 100 18788 400 18900
rect 100 18452 400 18564
rect 59600 18452 59900 18564
rect 100 17780 400 17892
rect 59600 17780 59900 17892
rect 59600 17444 59900 17556
rect 100 17108 400 17220
rect 100 16772 400 16884
rect 59600 16772 59900 16884
rect 100 16100 400 16212
rect 59600 16100 59900 16212
rect 59600 15764 59900 15876
rect 100 15428 400 15540
rect 59600 15092 59900 15204
rect 100 14756 400 14868
rect 100 14420 400 14532
rect 59600 14420 59900 14532
rect 100 13748 400 13860
rect 59600 13748 59900 13860
rect 59600 13412 59900 13524
rect 100 13076 400 13188
rect 59600 12740 59900 12852
rect 100 12404 400 12516
rect 100 12068 400 12180
rect 59600 12068 59900 12180
rect 100 11396 400 11508
rect 59600 11396 59900 11508
rect 59600 11060 59900 11172
rect 100 10724 400 10836
rect 100 10388 400 10500
rect 59600 10388 59900 10500
rect 100 9716 400 9828
rect 59600 9716 59900 9828
rect 59600 9380 59900 9492
rect 100 9044 400 9156
rect 59600 8708 59900 8820
rect 100 8372 400 8484
rect 100 8036 400 8148
rect 59600 8036 59900 8148
rect 100 7364 400 7476
rect 59600 7364 59900 7476
rect 59600 7028 59900 7140
rect 100 6692 400 6804
rect 59600 6356 59900 6468
rect 100 6020 400 6132
rect 100 5684 400 5796
rect 59600 5684 59900 5796
rect 100 5012 400 5124
rect 59600 5012 59900 5124
rect 59600 4676 59900 4788
rect 100 4340 400 4452
rect 100 4004 400 4116
rect 59600 4004 59900 4116
rect 100 3332 400 3444
rect 59600 3332 59900 3444
rect 59600 2996 59900 3108
rect 100 2660 400 2772
rect 59600 2324 59900 2436
rect 100 1988 400 2100
rect 100 1652 400 1764
rect 59600 1652 59900 1764
rect 100 980 400 1092
rect 59600 980 59900 1092
rect 59600 644 59900 756
rect 100 308 400 420
rect 59600 -28 59900 84
<< obsm3 >>
rect 65 59414 70 59458
rect 430 59414 59682 59458
rect 65 59250 59682 59414
rect 65 59078 59570 59250
rect 65 58914 59682 59078
rect 65 58742 70 58914
rect 430 58742 59682 58914
rect 65 58578 59682 58742
rect 65 58406 70 58578
rect 430 58406 59570 58578
rect 65 57906 59682 58406
rect 65 57734 70 57906
rect 430 57734 59570 57906
rect 65 57570 59682 57734
rect 65 57398 59570 57570
rect 65 57234 59682 57398
rect 65 57062 70 57234
rect 430 57062 59682 57234
rect 65 56898 59682 57062
rect 65 56726 70 56898
rect 430 56726 59570 56898
rect 65 56226 59682 56726
rect 65 56054 70 56226
rect 430 56054 59570 56226
rect 65 55890 59682 56054
rect 65 55718 59570 55890
rect 65 55554 59682 55718
rect 65 55382 70 55554
rect 430 55382 59682 55554
rect 65 55218 59682 55382
rect 65 55046 59570 55218
rect 65 54882 59682 55046
rect 65 54710 70 54882
rect 430 54710 59682 54882
rect 65 54546 59682 54710
rect 65 54374 70 54546
rect 430 54374 59570 54546
rect 65 53874 59682 54374
rect 65 53702 70 53874
rect 430 53702 59570 53874
rect 65 53538 59682 53702
rect 65 53366 59570 53538
rect 65 53202 59682 53366
rect 65 53030 70 53202
rect 430 53030 59682 53202
rect 65 52866 59682 53030
rect 65 52694 70 52866
rect 430 52694 59570 52866
rect 65 52194 59682 52694
rect 65 52022 70 52194
rect 430 52022 59570 52194
rect 65 51522 59682 52022
rect 65 51350 70 51522
rect 430 51350 59570 51522
rect 65 51186 59682 51350
rect 65 51014 59570 51186
rect 65 50850 59682 51014
rect 65 50678 70 50850
rect 430 50678 59682 50850
rect 65 50514 59682 50678
rect 65 50342 70 50514
rect 430 50342 59570 50514
rect 65 49842 59682 50342
rect 65 49670 70 49842
rect 430 49670 59570 49842
rect 65 49506 59682 49670
rect 65 49334 59570 49506
rect 65 49170 59682 49334
rect 65 48998 70 49170
rect 430 48998 59682 49170
rect 65 48834 59682 48998
rect 65 48662 59570 48834
rect 65 48498 59682 48662
rect 65 48326 70 48498
rect 430 48326 59682 48498
rect 65 48162 59682 48326
rect 65 47990 70 48162
rect 430 47990 59570 48162
rect 65 47490 59682 47990
rect 65 47318 70 47490
rect 430 47318 59570 47490
rect 65 47154 59682 47318
rect 65 46982 59570 47154
rect 65 46818 59682 46982
rect 65 46646 70 46818
rect 430 46646 59682 46818
rect 65 46482 59682 46646
rect 65 46310 70 46482
rect 430 46310 59570 46482
rect 65 45810 59682 46310
rect 65 45638 70 45810
rect 430 45638 59570 45810
rect 65 45474 59682 45638
rect 65 45302 59570 45474
rect 65 45138 59682 45302
rect 65 44966 70 45138
rect 430 44966 59682 45138
rect 65 44802 59682 44966
rect 65 44630 59570 44802
rect 65 44466 59682 44630
rect 65 44294 70 44466
rect 430 44294 59682 44466
rect 65 44130 59682 44294
rect 65 43958 70 44130
rect 430 43958 59570 44130
rect 65 43458 59682 43958
rect 65 43286 70 43458
rect 430 43286 59570 43458
rect 65 43122 59682 43286
rect 65 42950 59570 43122
rect 65 42786 59682 42950
rect 65 42614 70 42786
rect 430 42614 59682 42786
rect 65 42450 59682 42614
rect 65 42278 59570 42450
rect 65 42114 59682 42278
rect 65 41942 70 42114
rect 430 41942 59682 42114
rect 65 41778 59682 41942
rect 65 41606 70 41778
rect 430 41606 59570 41778
rect 65 41106 59682 41606
rect 65 40934 70 41106
rect 430 40934 59570 41106
rect 65 40770 59682 40934
rect 65 40598 59570 40770
rect 65 40434 59682 40598
rect 65 40262 70 40434
rect 430 40262 59682 40434
rect 65 40098 59682 40262
rect 65 39926 70 40098
rect 430 39926 59570 40098
rect 65 39426 59682 39926
rect 65 39254 70 39426
rect 430 39254 59570 39426
rect 65 39090 59682 39254
rect 65 38918 59570 39090
rect 65 38754 59682 38918
rect 65 38582 70 38754
rect 430 38582 59682 38754
rect 65 38418 59682 38582
rect 65 38246 59570 38418
rect 65 38082 59682 38246
rect 65 37910 70 38082
rect 430 37910 59682 38082
rect 65 37746 59682 37910
rect 65 37574 70 37746
rect 430 37574 59570 37746
rect 65 37074 59682 37574
rect 65 36902 70 37074
rect 430 36902 59570 37074
rect 65 36738 59682 36902
rect 65 36566 59570 36738
rect 65 36402 59682 36566
rect 65 36230 70 36402
rect 430 36230 59682 36402
rect 65 36066 59682 36230
rect 65 35894 59570 36066
rect 65 35730 59682 35894
rect 65 35558 70 35730
rect 430 35558 59682 35730
rect 65 35394 59682 35558
rect 65 35222 70 35394
rect 430 35222 59570 35394
rect 65 34722 59682 35222
rect 65 34550 70 34722
rect 430 34550 59570 34722
rect 65 34386 59682 34550
rect 65 34214 59570 34386
rect 65 34050 59682 34214
rect 65 33878 70 34050
rect 430 33878 59682 34050
rect 65 33714 59682 33878
rect 65 33542 70 33714
rect 430 33542 59570 33714
rect 65 33042 59682 33542
rect 65 32870 70 33042
rect 430 32870 59570 33042
rect 65 32706 59682 32870
rect 65 32534 59570 32706
rect 65 32370 59682 32534
rect 65 32198 70 32370
rect 430 32198 59682 32370
rect 65 32034 59682 32198
rect 65 31862 59570 32034
rect 65 31698 59682 31862
rect 65 31526 70 31698
rect 430 31526 59682 31698
rect 65 31362 59682 31526
rect 65 31190 70 31362
rect 430 31190 59570 31362
rect 65 30690 59682 31190
rect 65 30518 70 30690
rect 430 30518 59570 30690
rect 65 30354 59682 30518
rect 65 30182 59570 30354
rect 65 30018 59682 30182
rect 65 29846 70 30018
rect 430 29846 59682 30018
rect 65 29682 59682 29846
rect 65 29510 59570 29682
rect 65 29346 59682 29510
rect 65 29174 70 29346
rect 430 29174 59682 29346
rect 65 29010 59682 29174
rect 65 28838 70 29010
rect 430 28838 59570 29010
rect 65 28338 59682 28838
rect 65 28166 70 28338
rect 430 28166 59570 28338
rect 65 28002 59682 28166
rect 65 27830 59570 28002
rect 65 27666 59682 27830
rect 65 27494 70 27666
rect 430 27494 59682 27666
rect 65 27330 59682 27494
rect 65 27158 70 27330
rect 430 27158 59570 27330
rect 65 26658 59682 27158
rect 65 26486 70 26658
rect 430 26486 59570 26658
rect 65 26322 59682 26486
rect 65 26150 59570 26322
rect 65 25986 59682 26150
rect 65 25814 70 25986
rect 430 25814 59682 25986
rect 65 25650 59682 25814
rect 65 25478 59570 25650
rect 65 25314 59682 25478
rect 65 25142 70 25314
rect 430 25142 59682 25314
rect 65 24978 59682 25142
rect 65 24806 70 24978
rect 430 24806 59570 24978
rect 65 24306 59682 24806
rect 65 24134 70 24306
rect 430 24134 59570 24306
rect 65 23970 59682 24134
rect 65 23798 59570 23970
rect 65 23634 59682 23798
rect 65 23462 70 23634
rect 430 23462 59682 23634
rect 65 23298 59682 23462
rect 65 23126 70 23298
rect 430 23126 59570 23298
rect 65 22626 59682 23126
rect 65 22454 70 22626
rect 430 22454 59570 22626
rect 65 21954 59682 22454
rect 65 21782 70 21954
rect 430 21782 59570 21954
rect 65 21618 59682 21782
rect 65 21446 59570 21618
rect 65 21282 59682 21446
rect 65 21110 70 21282
rect 430 21110 59682 21282
rect 65 20946 59682 21110
rect 65 20774 70 20946
rect 430 20774 59570 20946
rect 65 20274 59682 20774
rect 65 20102 70 20274
rect 430 20102 59570 20274
rect 65 19938 59682 20102
rect 65 19766 59570 19938
rect 65 19602 59682 19766
rect 65 19430 70 19602
rect 430 19430 59682 19602
rect 65 19266 59682 19430
rect 65 19094 59570 19266
rect 65 18930 59682 19094
rect 65 18758 70 18930
rect 430 18758 59682 18930
rect 65 18594 59682 18758
rect 65 18422 70 18594
rect 430 18422 59570 18594
rect 65 17922 59682 18422
rect 65 17750 70 17922
rect 430 17750 59570 17922
rect 65 17586 59682 17750
rect 65 17414 59570 17586
rect 65 17250 59682 17414
rect 65 17078 70 17250
rect 430 17078 59682 17250
rect 65 16914 59682 17078
rect 65 16742 70 16914
rect 430 16742 59570 16914
rect 65 16242 59682 16742
rect 65 16070 70 16242
rect 430 16070 59570 16242
rect 65 15906 59682 16070
rect 65 15734 59570 15906
rect 65 15570 59682 15734
rect 65 15398 70 15570
rect 430 15398 59682 15570
rect 65 15234 59682 15398
rect 65 15062 59570 15234
rect 65 14898 59682 15062
rect 65 14726 70 14898
rect 430 14726 59682 14898
rect 65 14562 59682 14726
rect 65 14390 70 14562
rect 430 14390 59570 14562
rect 65 13890 59682 14390
rect 65 13718 70 13890
rect 430 13718 59570 13890
rect 65 13554 59682 13718
rect 65 13382 59570 13554
rect 65 13218 59682 13382
rect 65 13046 70 13218
rect 430 13046 59682 13218
rect 65 12882 59682 13046
rect 65 12710 59570 12882
rect 65 12546 59682 12710
rect 65 12374 70 12546
rect 430 12374 59682 12546
rect 65 12210 59682 12374
rect 65 12038 70 12210
rect 430 12038 59570 12210
rect 65 11538 59682 12038
rect 65 11366 70 11538
rect 430 11366 59570 11538
rect 65 11202 59682 11366
rect 65 11030 59570 11202
rect 65 10866 59682 11030
rect 65 10694 70 10866
rect 430 10694 59682 10866
rect 65 10530 59682 10694
rect 65 10358 70 10530
rect 430 10358 59570 10530
rect 65 9858 59682 10358
rect 65 9686 70 9858
rect 430 9686 59570 9858
rect 65 9522 59682 9686
rect 65 9350 59570 9522
rect 65 9186 59682 9350
rect 65 9014 70 9186
rect 430 9014 59682 9186
rect 65 8850 59682 9014
rect 65 8678 59570 8850
rect 65 8514 59682 8678
rect 65 8342 70 8514
rect 430 8342 59682 8514
rect 65 8178 59682 8342
rect 65 8006 70 8178
rect 430 8006 59570 8178
rect 65 7506 59682 8006
rect 65 7334 70 7506
rect 430 7334 59570 7506
rect 65 7170 59682 7334
rect 65 6998 59570 7170
rect 65 6834 59682 6998
rect 65 6662 70 6834
rect 430 6662 59682 6834
rect 65 6498 59682 6662
rect 65 6326 59570 6498
rect 65 6162 59682 6326
rect 65 5990 70 6162
rect 430 5990 59682 6162
rect 65 5826 59682 5990
rect 65 5654 70 5826
rect 430 5654 59570 5826
rect 65 5154 59682 5654
rect 65 4982 70 5154
rect 430 4982 59570 5154
rect 65 4818 59682 4982
rect 65 4646 59570 4818
rect 65 4482 59682 4646
rect 65 4310 70 4482
rect 430 4310 59682 4482
rect 65 4146 59682 4310
rect 65 3974 70 4146
rect 430 3974 59570 4146
rect 65 3474 59682 3974
rect 65 3302 70 3474
rect 430 3302 59570 3474
rect 65 3138 59682 3302
rect 65 2966 59570 3138
rect 65 2802 59682 2966
rect 65 2630 70 2802
rect 430 2630 59682 2802
rect 65 2466 59682 2630
rect 65 2294 59570 2466
rect 65 2130 59682 2294
rect 65 1958 70 2130
rect 430 1958 59682 2130
rect 65 1794 59682 1958
rect 65 1622 70 1794
rect 430 1622 59570 1794
rect 65 1122 59682 1622
rect 65 950 70 1122
rect 430 950 59570 1122
rect 65 786 59682 950
rect 65 742 59570 786
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 23870 21849 25234 31687
rect 25454 21849 32914 31687
rect 33134 21849 36666 31687
<< labels >>
rlabel metal3 s 100 20804 400 20916 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 27524 400 27636 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 24836 400 24948 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57764 59600 57876 59900 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 21140 400 21252 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 32900 59600 33012 59900 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 59600 11396 59900 11508 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 17108 100 17220 400 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 13412 59600 13524 59900 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 26516 400 26628 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 59600 59780 59900 59892 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 48020 59600 48132 59900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 34580 59600 34692 59900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 56756 59600 56868 59900 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 980 59600 1092 59900 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 8036 100 8148 400 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 7364 59600 7476 59900 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 9716 59600 9828 59900 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 59600 6356 59900 6468 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 14420 400 14532 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 2324 59600 2436 59900 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 59600 58436 59900 58548 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 6020 400 6132 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 41972 100 42084 400 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 8708 59600 8820 59900 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 35588 100 35700 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 58772 400 58884 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53732 59600 53844 59900 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 12740 59600 12852 59900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 100 15428 400 15540 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59600 9716 59900 9828 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 25172 400 25284 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 53732 100 53844 400 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 58436 400 58548 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 100 13748 400 13860 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 59600 15764 59900 15876 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 58436 100 58548 400 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 51044 59600 51156 59900 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1652 59600 1764 59900 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 100 40964 400 41076 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 37604 400 37716 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 100 44996 400 45108 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 51380 100 51492 400 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 58772 100 58884 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 31892 59600 32004 59900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 100 34580 400 34692 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 5684 59600 5796 59900 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 47348 400 47460 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 24164 100 24276 400 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 59600 4676 59900 4788 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 50708 100 50820 400 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 5684 100 5796 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 59600 15092 59900 15204 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 100 5684 400 5796 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 59600 13412 59900 13524 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 21140 100 21252 400 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 49700 100 49812 400 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 100 39956 400 40068 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 56084 400 56196 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 12068 59600 12180 59900 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 38612 100 38724 400 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 100 1988 400 2100 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 59600 41636 59900 41748 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 59600 9380 59900 9492 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 100 49028 400 49140 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 23156 400 23268 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 33572 59600 33684 59900 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 56084 100 56196 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 50372 400 50484 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 59600 20132 59900 20244 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s -28 59600 84 59900 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 59600 57764 59900 57876 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 28868 59600 28980 59900 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 59600 3332 59900 3444 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 59600 24164 59900 24276 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 59600 23828 59900 23940 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 100 11396 400 11508 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 58436 59600 58548 59900 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 59600 52724 59900 52836 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 59600 59108 59900 59220 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 44324 400 44436 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23492 100 23604 400 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 59600 49700 59900 49812 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 6692 100 6804 400 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 50372 100 50484 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 39284 100 39396 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 4004 100 4116 400 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 40964 100 41076 400 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 27188 100 27300 400 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 20132 100 20244 400 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 100 8036 400 8148 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 43988 59600 44100 59900 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 27860 59600 27972 59900 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 25172 100 25284 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42308 59600 42420 59900 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 44324 100 44436 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 38276 59600 38388 59900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 56756 100 56868 400 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 55076 59600 55188 59900 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 59600 12740 59900 12852 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50372 59600 50484 59900 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 59600 19124 59900 19236 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 39956 100 40068 400 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 59600 38948 59900 39060 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 14420 100 14532 400 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 59600 56084 59900 56196 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 59600 55748 59900 55860 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 59600 42980 59900 43092 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 100 1652 400 1764 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 100 2660 400 2772 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 33908 400 34020 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37604 59600 37716 59900 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 15428 100 15540 400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 30548 400 30660 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 41972 400 42084 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 100 24164 400 24276 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 18452 100 18564 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 24164 59600 24276 59900 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 56084 59600 56196 59900 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 28196 100 28308 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal3 s 100 36260 400 36372 6 la_data_in[12]
port 121 nsew signal input
rlabel metal3 s 59600 8708 59900 8820 6 la_data_in[13]
port 122 nsew signal input
rlabel metal3 s 59600 21812 59900 21924 6 la_data_in[14]
port 123 nsew signal input
rlabel metal3 s 100 41636 400 41748 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 13748 59600 13860 59900 6 la_data_in[16]
port 125 nsew signal input
rlabel metal3 s 59600 12068 59900 12180 6 la_data_in[17]
port 126 nsew signal input
rlabel metal3 s 59600 45332 59900 45444 6 la_data_in[18]
port 127 nsew signal input
rlabel metal3 s 59600 26516 59900 26628 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 45668 59600 45780 59900 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 30548 59600 30660 59900 6 la_data_in[20]
port 130 nsew signal input
rlabel metal3 s 100 9716 400 9828 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 36932 59600 37044 59900 6 la_data_in[22]
port 132 nsew signal input
rlabel metal3 s 100 54404 400 54516 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 26180 59600 26292 59900 6 la_data_in[24]
port 134 nsew signal input
rlabel metal3 s 59600 14420 59900 14532 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 19460 100 19572 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal3 s 100 4340 400 4452 6 la_data_in[27]
port 137 nsew signal input
rlabel metal3 s 100 21812 400 21924 6 la_data_in[28]
port 138 nsew signal input
rlabel metal3 s 100 45668 400 45780 6 la_data_in[29]
port 139 nsew signal input
rlabel metal3 s 100 40292 400 40404 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 4676 59600 4788 59900 6 la_data_in[30]
port 141 nsew signal input
rlabel metal3 s 100 53060 400 53172 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 30212 59600 30324 59900 6 la_data_in[32]
port 143 nsew signal input
rlabel metal3 s 59600 51044 59900 51156 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 18452 59600 18564 59900 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 24836 59600 24948 59900 6 la_data_in[35]
port 146 nsew signal input
rlabel metal3 s 59600 32564 59900 32676 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 20804 100 20916 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 28868 100 28980 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal3 s 100 20132 400 20244 6 la_data_in[39]
port 150 nsew signal input
rlabel metal3 s 59600 36932 59900 37044 6 la_data_in[3]
port 151 nsew signal input
rlabel metal3 s 59600 644 59900 756 6 la_data_in[40]
port 152 nsew signal input
rlabel metal3 s 100 56756 400 56868 6 la_data_in[41]
port 153 nsew signal input
rlabel metal3 s 59600 43316 59900 43428 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 36932 100 37044 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 28196 59600 28308 59900 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 8036 59600 8148 59900 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 5012 59600 5124 59900 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 23828 59600 23940 59900 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 27524 100 27636 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal3 s 100 31220 400 31332 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 49364 59600 49476 59900 6 la_data_in[4]
port 162 nsew signal input
rlabel metal3 s 100 18452 400 18564 6 la_data_in[50]
port 163 nsew signal input
rlabel metal3 s 100 16100 400 16212 6 la_data_in[51]
port 164 nsew signal input
rlabel metal3 s 100 17780 400 17892 6 la_data_in[52]
port 165 nsew signal input
rlabel metal3 s 59600 1652 59900 1764 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 21812 100 21924 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal3 s 59600 54404 59900 54516 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 10388 100 10500 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 15764 59600 15876 59900 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 22484 59600 22596 59900 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 35252 100 35364 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal3 s 100 308 400 420 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 12068 100 12180 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal3 s 59600 21476 59900 21588 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 17780 59600 17892 59900 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 54404 59600 54516 59900 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 52052 59600 52164 59900 6 la_data_in[6]
port 178 nsew signal input
rlabel metal3 s 59600 31892 59900 32004 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 42644 100 42756 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal3 s 100 43316 400 43428 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 16772 59600 16884 59900 6 la_data_out[0]
port 182 nsew signal output
rlabel metal3 s 59600 24836 59900 24948 6 la_data_out[10]
port 183 nsew signal output
rlabel metal3 s 100 51380 400 51492 6 la_data_out[11]
port 184 nsew signal output
rlabel metal3 s 59600 32900 59900 33012 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 29540 59600 29652 59900 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 26516 59600 26628 59900 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 31556 100 31668 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal3 s 59600 27860 59900 27972 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 59108 59600 59220 59900 6 la_data_out[17]
port 190 nsew signal output
rlabel metal3 s 100 59444 400 59556 6 la_data_out[18]
port 191 nsew signal output
rlabel metal3 s 59600 37604 59900 37716 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 17780 100 17892 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal3 s 59600 17444 59900 17556 6 la_data_out[20]
port 194 nsew signal output
rlabel metal3 s 100 10388 400 10500 6 la_data_out[21]
port 195 nsew signal output
rlabel metal3 s 59600 7364 59900 7476 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 36596 59600 36708 59900 6 la_data_out[23]
port 197 nsew signal output
rlabel metal3 s 59600 47348 59900 47460 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 25844 100 25956 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal3 s 100 46676 400 46788 6 la_data_out[26]
port 200 nsew signal output
rlabel metal3 s 59600 27188 59900 27300 6 la_data_out[27]
port 201 nsew signal output
rlabel metal3 s 100 22484 400 22596 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 35252 59600 35364 59900 6 la_data_out[29]
port 203 nsew signal output
rlabel metal3 s 59600 11060 59900 11172 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 29204 100 29316 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 32564 59600 32676 59900 6 la_data_out[31]
port 206 nsew signal output
rlabel metal3 s 59600 48020 59900 48132 6 la_data_out[32]
port 207 nsew signal output
rlabel metal3 s 59600 23156 59900 23268 6 la_data_out[33]
port 208 nsew signal output
rlabel metal3 s 59600 980 59900 1092 6 la_data_out[34]
port 209 nsew signal output
rlabel metal3 s 59600 8036 59900 8148 6 la_data_out[35]
port 210 nsew signal output
rlabel metal3 s 100 3332 400 3444 6 la_data_out[36]
port 211 nsew signal output
rlabel metal3 s 100 53732 400 53844 6 la_data_out[37]
port 212 nsew signal output
rlabel metal3 s 100 27188 400 27300 6 la_data_out[38]
port 213 nsew signal output
rlabel metal3 s 59600 50372 59900 50484 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 3332 100 3444 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 24836 100 24948 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 9380 59600 9492 59900 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 54740 100 54852 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal3 s 100 42644 400 42756 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 13748 100 13860 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 54404 100 54516 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 34244 59600 34356 59900 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 20804 59600 20916 59900 6 la_data_out[47]
port 223 nsew signal output
rlabel metal3 s 100 57764 400 57876 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 43316 59600 43428 59900 6 la_data_out[49]
port 225 nsew signal output
rlabel metal3 s 100 980 400 1092 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 47012 59600 47124 59900 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 25508 59600 25620 59900 6 la_data_out[51]
port 228 nsew signal output
rlabel metal3 s 100 8372 400 8484 6 la_data_out[52]
port 229 nsew signal output
rlabel metal3 s 59600 35252 59900 35364 6 la_data_out[53]
port 230 nsew signal output
rlabel metal3 s 59600 40964 59900 41076 6 la_data_out[54]
port 231 nsew signal output
rlabel metal3 s 59600 53396 59900 53508 6 la_data_out[55]
port 232 nsew signal output
rlabel metal3 s 100 54740 400 54852 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 48692 59600 48804 59900 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 16100 100 16212 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 52052 100 52164 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal3 s 59600 4004 59900 4116 6 la_data_out[5]
port 237 nsew signal output
rlabel metal3 s 100 9044 400 9156 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 21476 59600 21588 59900 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 37604 100 37716 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal3 s 59600 28196 59900 28308 6 la_data_out[63]
port 241 nsew signal output
rlabel metal3 s 59600 22484 59900 22596 6 la_data_out[6]
port 242 nsew signal output
rlabel metal3 s 59600 42308 59900 42420 6 la_data_out[7]
port 243 nsew signal output
rlabel metal3 s 59600 33572 59900 33684 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 23156 59600 23268 59900 6 la_data_out[9]
port 245 nsew signal output
rlabel metal3 s 100 48020 400 48132 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 43988 100 44100 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 52724 100 52836 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 8372 100 8484 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal3 s 100 7364 400 7476 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 4004 59600 4116 59900 6 la_oenb[14]
port 251 nsew signal input
rlabel metal3 s 59600 5012 59900 5124 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 11396 59600 11508 59900 6 la_oenb[16]
port 253 nsew signal input
rlabel metal3 s 100 52724 400 52836 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 52724 59600 52836 59900 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 44660 59600 44772 59900 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 16772 100 16884 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal3 s 100 33572 400 33684 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 53060 100 53172 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal3 s 100 32228 400 32340 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 10724 100 10836 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal3 s 100 36932 400 37044 6 la_oenb[24]
port 262 nsew signal input
rlabel metal3 s 59600 56756 59900 56868 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 59780 59600 59892 59900 6 la_oenb[26]
port 264 nsew signal input
rlabel metal3 s 59600 51380 59900 51492 6 la_oenb[27]
port 265 nsew signal input
rlabel metal3 s 59600 49364 59900 49476 6 la_oenb[28]
port 266 nsew signal input
rlabel metal3 s 59600 48692 59900 48804 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 30548 100 30660 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 10388 59600 10500 59900 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 1652 100 1764 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 308 100 420 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 644 59600 756 59900 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 31220 100 31332 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal3 s 100 25844 400 25956 6 la_oenb[35]
port 274 nsew signal input
rlabel metal3 s 100 32900 400 33012 6 la_oenb[36]
port 275 nsew signal input
rlabel metal3 s 100 17108 400 17220 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 21812 59600 21924 59900 6 la_oenb[38]
port 277 nsew signal input
rlabel metal3 s 100 37940 400 38052 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 11396 100 11508 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 26516 100 26628 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal3 s 100 29876 400 29988 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 48020 100 48132 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 22484 100 22596 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal3 s 100 43988 400 44100 6 la_oenb[44]
port 284 nsew signal input
rlabel metal3 s 59600 28868 59900 28980 6 la_oenb[45]
port 285 nsew signal input
rlabel metal3 s 59600 39956 59900 40068 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 46340 100 46452 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 19796 59600 19908 59900 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 59444 100 59556 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal3 s 59600 38276 59900 38388 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 40628 59600 40740 59900 6 la_oenb[50]
port 291 nsew signal input
rlabel metal3 s 59600 30548 59900 30660 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 45668 100 45780 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 53396 59600 53508 59900 6 la_oenb[53]
port 294 nsew signal input
rlabel metal3 s 59600 5684 59900 5796 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 35924 59600 36036 59900 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 55412 100 55524 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal3 s 100 29204 400 29316 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 7364 100 7476 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal3 s 59600 30212 59900 30324 6 la_oenb[59]
port 300 nsew signal input
rlabel metal3 s 100 57092 400 57204 6 la_oenb[5]
port 301 nsew signal input
rlabel metal3 s 59600 39284 59900 39396 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 14756 100 14868 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 57092 100 57204 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal3 s 100 10724 400 10836 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 51380 59600 51492 59900 6 la_oenb[6]
port 306 nsew signal input
rlabel metal3 s 59600 45668 59900 45780 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 15092 59600 15204 59900 6 la_oenb[8]
port 308 nsew signal input
rlabel metal3 s 100 38612 400 38724 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal3 s 59600 10388 59900 10500 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 11060 59600 11172 59900 6 wb_rst_i
port 313 nsew signal input
rlabel metal3 s 59600 20804 59900 20916 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 39956 59600 40068 59900 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 27188 59600 27300 59900 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 3332 59600 3444 59900 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 5012 100 5124 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 33572 100 33684 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal3 s 59600 43988 59900 44100 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal3 s 59600 40628 59900 40740 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 37940 100 38052 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal3 s 59600 35924 59900 36036 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal3 s 59600 18452 59900 18564 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 57764 100 57876 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal3 s 100 4004 400 4116 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal3 s 100 35252 400 35364 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 33908 100 34020 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 48356 100 48468 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal3 s 59600 13748 59900 13860 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 7028 59600 7140 59900 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 32900 100 33012 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 6020 100 6132 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 20132 59600 20244 59900 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal3 s 59600 34580 59900 34692 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal3 s 59600 57428 59900 57540 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal3 s 100 6692 400 6804 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal3 s 100 23492 400 23604 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal3 s 59600 25508 59900 25620 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 46676 100 46788 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 46340 59600 46452 59900 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 44996 100 45108 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal3 s 100 28868 400 28980 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 2660 100 2772 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal3 s 59600 -28 59900 84 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal3 s 59600 16100 59900 16212 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 19124 59600 19236 59900 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal3 s 59600 52052 59900 52164 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal3 s 100 46340 400 46452 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal3 s 100 50708 400 50820 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal3 s 100 48356 400 48468 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 1988 100 2100 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal3 s 100 12404 400 12516 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal3 s 59600 31220 59900 31332 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 34580 100 34692 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 40964 59600 41076 59900 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 55748 59600 55860 59900 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 2996 59600 3108 59900 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 9044 100 9156 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal3 s 100 14756 400 14868 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 57428 59600 57540 59900 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal3 s 100 35588 400 35700 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal3 s 59600 47012 59900 47124 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal3 s 59600 19796 59900 19908 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 41636 100 41748 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 49700 59600 49812 59900 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 14420 59600 14532 59900 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 18788 100 18900 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal3 s 59600 36596 59900 36708 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 49028 100 49140 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal3 s 59600 17780 59900 17892 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal3 s 100 31556 400 31668 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal3 s 59600 2324 59900 2436 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 9716 100 9828 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 29876 100 29988 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal3 s 59600 26180 59900 26292 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 47348 59600 47460 59900 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal3 s 59600 53732 59900 53844 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal3 s 59600 2996 59900 3108 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal3 s 100 12068 400 12180 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal3 s 59600 34244 59900 34356 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 980 100 1092 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal3 s 59600 55076 59900 55188 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 45332 59600 45444 59900 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal3 s 59600 7028 59900 7140 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 42980 59600 43092 59900 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal3 s 100 16772 400 16884 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal3 s 100 18788 400 18900 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 40292 100 40404 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s -28 100 84 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 47348 100 47460 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal3 s 100 28196 400 28308 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal3 s 100 52052 400 52164 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 16100 59600 16212 59900 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal3 s 100 19460 400 19572 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 12404 100 12516 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 4340 100 4452 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 31220 59600 31332 59900 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 17444 59600 17556 59900 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 32228 100 32340 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 41636 59600 41748 59900 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal3 s 59600 16772 59900 16884 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal3 s 100 39284 400 39396 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal3 s 59600 46340 59900 46452 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 13076 100 13188 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 23156 100 23268 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal3 s 100 5012 400 5124 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal3 s 59600 44660 59900 44772 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 36260 100 36372 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 39284 59600 39396 59900 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 38948 59600 39060 59900 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal3 s 100 55412 400 55524 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 6356 59600 6468 59900 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 43316 100 43428 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal3 s 100 13076 400 13188 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal3 s 100 49700 400 49812 6 wbs_stb_i
port 416 nsew signal input
rlabel metal3 s 59600 29540 59900 29652 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2886700
string GDS_FILE /home/dastechlabs/FPGA_Projects/Fuzzy-Wavelet_Clone/caravel_user_project/openlane/wrapped_fuzzy_wavelet/runs/22_12_05_16_37/results/signoff/user_proj_example.magic.gds
string GDS_START 238166
<< end >>

