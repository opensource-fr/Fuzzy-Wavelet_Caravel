magic
tech gf180mcuC
magscale 1 10
timestamp 1670287216
<< metal1 >>
rect 1698 117070 1710 117122
rect 1762 117119 1774 117122
rect 1922 117119 1934 117122
rect 1762 117073 1934 117119
rect 1762 117070 1774 117073
rect 1922 117070 1934 117073
rect 1986 117070 1998 117122
rect 39778 117070 39790 117122
rect 39842 117119 39854 117122
rect 41122 117119 41134 117122
rect 39842 117073 41134 117119
rect 39842 117070 39854 117073
rect 41122 117070 41134 117073
rect 41186 117070 41198 117122
rect 63970 116958 63982 117010
rect 64034 117007 64046 117010
rect 65202 117007 65214 117010
rect 64034 116961 65214 117007
rect 64034 116958 64046 116961
rect 65202 116958 65214 116961
rect 65266 116958 65278 117010
rect 67218 116958 67230 117010
rect 67282 117007 67294 117010
rect 68450 117007 68462 117010
rect 67282 116961 68462 117007
rect 67282 116958 67294 116961
rect 68450 116958 68462 116961
rect 68514 116958 68526 117010
rect 1344 116842 118608 116876
rect 1344 116790 4478 116842
rect 4530 116790 4582 116842
rect 4634 116790 4686 116842
rect 4738 116790 35198 116842
rect 35250 116790 35302 116842
rect 35354 116790 35406 116842
rect 35458 116790 65918 116842
rect 65970 116790 66022 116842
rect 66074 116790 66126 116842
rect 66178 116790 96638 116842
rect 96690 116790 96742 116842
rect 96794 116790 96846 116842
rect 96898 116790 118608 116842
rect 1344 116756 118608 116790
rect 5854 116562 5906 116574
rect 9886 116562 9938 116574
rect 12798 116562 12850 116574
rect 21982 116562 22034 116574
rect 36990 116562 37042 116574
rect 3266 116510 3278 116562
rect 3330 116510 3342 116562
rect 7522 116510 7534 116562
rect 7586 116510 7598 116562
rect 11778 116510 11790 116562
rect 11842 116510 11854 116562
rect 16706 116510 16718 116562
rect 16770 116510 16782 116562
rect 23874 116510 23886 116562
rect 23938 116510 23950 116562
rect 26002 116510 26014 116562
rect 26066 116510 26078 116562
rect 32162 116510 32174 116562
rect 32226 116510 32238 116562
rect 36306 116510 36318 116562
rect 36370 116510 36382 116562
rect 5854 116498 5906 116510
rect 9886 116498 9938 116510
rect 12798 116498 12850 116510
rect 21982 116498 22034 116510
rect 36990 116498 37042 116510
rect 37438 116562 37490 116574
rect 37438 116498 37490 116510
rect 38110 116562 38162 116574
rect 45054 116562 45106 116574
rect 49534 116562 49586 116574
rect 56030 116562 56082 116574
rect 59950 116562 60002 116574
rect 81118 116562 81170 116574
rect 95118 116562 95170 116574
rect 99150 116562 99202 116574
rect 106878 116562 106930 116574
rect 110910 116562 110962 116574
rect 114830 116562 114882 116574
rect 39778 116510 39790 116562
rect 39842 116510 39854 116562
rect 48066 116510 48078 116562
rect 48130 116510 48142 116562
rect 51202 116510 51214 116562
rect 51266 116510 51278 116562
rect 54002 116510 54014 116562
rect 54066 116510 54078 116562
rect 58146 116510 58158 116562
rect 58210 116510 58222 116562
rect 60946 116510 60958 116562
rect 61010 116510 61022 116562
rect 65202 116510 65214 116562
rect 65266 116510 65278 116562
rect 66434 116510 66446 116562
rect 66498 116510 66510 116562
rect 69122 116510 69134 116562
rect 69186 116510 69198 116562
rect 70578 116510 70590 116562
rect 70642 116510 70654 116562
rect 72482 116510 72494 116562
rect 72546 116510 72558 116562
rect 76962 116510 76974 116562
rect 77026 116510 77038 116562
rect 78978 116510 78990 116562
rect 79042 116510 79054 116562
rect 81554 116510 81566 116562
rect 81618 116510 81630 116562
rect 84802 116510 84814 116562
rect 84866 116510 84878 116562
rect 86594 116510 86606 116562
rect 86658 116510 86670 116562
rect 89058 116510 89070 116562
rect 89122 116510 89134 116562
rect 92642 116510 92654 116562
rect 92706 116510 92718 116562
rect 95890 116510 95902 116562
rect 95954 116510 95966 116562
rect 99810 116510 99822 116562
rect 99874 116510 99886 116562
rect 107650 116510 107662 116562
rect 107714 116510 107726 116562
rect 111794 116510 111806 116562
rect 111858 116510 111870 116562
rect 115714 116510 115726 116562
rect 115778 116510 115790 116562
rect 38110 116498 38162 116510
rect 45054 116498 45106 116510
rect 49534 116498 49586 116510
rect 56030 116498 56082 116510
rect 59950 116498 60002 116510
rect 81118 116498 81170 116510
rect 95118 116498 95170 116510
rect 99150 116498 99202 116510
rect 106878 116498 106930 116510
rect 110910 116498 110962 116510
rect 114830 116498 114882 116510
rect 17390 116450 17442 116462
rect 4050 116398 4062 116450
rect 4114 116398 4126 116450
rect 25330 116398 25342 116450
rect 25394 116398 25406 116450
rect 53330 116398 53342 116450
rect 53394 116398 53406 116450
rect 64530 116398 64542 116450
rect 64594 116398 64606 116450
rect 67554 116398 67566 116450
rect 67618 116398 67630 116450
rect 68450 116398 68462 116450
rect 68514 116398 68526 116450
rect 71362 116398 71374 116450
rect 71426 116398 71438 116450
rect 76290 116398 76302 116450
rect 76354 116398 76366 116450
rect 78194 116398 78206 116450
rect 78258 116398 78270 116450
rect 84130 116398 84142 116450
rect 84194 116398 84206 116450
rect 85922 116398 85934 116450
rect 85986 116398 85998 116450
rect 88274 116398 88286 116450
rect 88338 116398 88350 116450
rect 91970 116398 91982 116450
rect 92034 116398 92046 116450
rect 17390 116386 17442 116398
rect 19070 116338 19122 116350
rect 33070 116338 33122 116350
rect 44046 116338 44098 116350
rect 48750 116338 48802 116350
rect 94334 116338 94386 116350
rect 97918 116338 97970 116350
rect 1922 116286 1934 116338
rect 1986 116286 1998 116338
rect 6402 116286 6414 116338
rect 6466 116286 6478 116338
rect 10434 116286 10446 116338
rect 10498 116286 10510 116338
rect 15698 116286 15710 116338
rect 15762 116286 15774 116338
rect 22530 116286 22542 116338
rect 22594 116286 22606 116338
rect 31378 116286 31390 116338
rect 31442 116286 31454 116338
rect 35186 116286 35198 116338
rect 35250 116286 35262 116338
rect 38658 116286 38670 116338
rect 38722 116286 38734 116338
rect 41122 116286 41134 116338
rect 41186 116286 41198 116338
rect 46946 116286 46958 116338
rect 47010 116286 47022 116338
rect 50082 116286 50094 116338
rect 50146 116286 50158 116338
rect 56802 116286 56814 116338
rect 56866 116286 56878 116338
rect 61730 116286 61742 116338
rect 61794 116286 61806 116338
rect 74386 116286 74398 116338
rect 74450 116286 74462 116338
rect 82562 116286 82574 116338
rect 82626 116286 82638 116338
rect 96898 116286 96910 116338
rect 96962 116286 96974 116338
rect 100818 116286 100830 116338
rect 100882 116286 100894 116338
rect 108658 116286 108670 116338
rect 108722 116286 108734 116338
rect 112802 116286 112814 116338
rect 112866 116286 112878 116338
rect 116498 116286 116510 116338
rect 116562 116286 116574 116338
rect 19070 116274 19122 116286
rect 33070 116274 33122 116286
rect 44046 116274 44098 116286
rect 48750 116274 48802 116286
rect 94334 116274 94386 116286
rect 97918 116274 97970 116286
rect 3838 116226 3890 116238
rect 3838 116162 3890 116174
rect 4734 116226 4786 116238
rect 4734 116162 4786 116174
rect 43598 116226 43650 116238
rect 43598 116162 43650 116174
rect 52782 116226 52834 116238
rect 52782 116162 52834 116174
rect 75518 116226 75570 116238
rect 75518 116162 75570 116174
rect 91198 116226 91250 116238
rect 91198 116162 91250 116174
rect 117518 116226 117570 116238
rect 117518 116162 117570 116174
rect 1344 116058 118608 116092
rect 1344 116006 19838 116058
rect 19890 116006 19942 116058
rect 19994 116006 20046 116058
rect 20098 116006 50558 116058
rect 50610 116006 50662 116058
rect 50714 116006 50766 116058
rect 50818 116006 81278 116058
rect 81330 116006 81382 116058
rect 81434 116006 81486 116058
rect 81538 116006 111998 116058
rect 112050 116006 112102 116058
rect 112154 116006 112206 116058
rect 112258 116006 118608 116058
rect 1344 115972 118608 116006
rect 5742 115890 5794 115902
rect 5742 115826 5794 115838
rect 22766 115890 22818 115902
rect 22766 115826 22818 115838
rect 23550 115890 23602 115902
rect 23550 115826 23602 115838
rect 24110 115890 24162 115902
rect 24110 115826 24162 115838
rect 28702 115890 28754 115902
rect 28702 115826 28754 115838
rect 40798 115890 40850 115902
rect 40798 115826 40850 115838
rect 41918 115890 41970 115902
rect 41918 115826 41970 115838
rect 51326 115890 51378 115902
rect 51326 115826 51378 115838
rect 67230 115890 67282 115902
rect 67230 115826 67282 115838
rect 68686 115890 68738 115902
rect 68686 115826 68738 115838
rect 69582 115890 69634 115902
rect 69582 115826 69634 115838
rect 81790 115890 81842 115902
rect 81790 115826 81842 115838
rect 85262 115890 85314 115902
rect 85262 115826 85314 115838
rect 108670 115890 108722 115902
rect 108670 115826 108722 115838
rect 10670 115778 10722 115790
rect 72606 115778 72658 115790
rect 1922 115726 1934 115778
rect 1986 115726 1998 115778
rect 3714 115726 3726 115778
rect 3778 115726 3790 115778
rect 13122 115726 13134 115778
rect 13186 115726 13198 115778
rect 29250 115726 29262 115778
rect 29314 115726 29326 115778
rect 35298 115726 35310 115778
rect 35362 115726 35374 115778
rect 37314 115726 37326 115778
rect 37378 115726 37390 115778
rect 43586 115726 43598 115778
rect 43650 115726 43662 115778
rect 45378 115726 45390 115778
rect 45442 115726 45454 115778
rect 62850 115726 62862 115778
rect 62914 115726 62926 115778
rect 78978 115726 78990 115778
rect 79042 115726 79054 115778
rect 83234 115726 83246 115778
rect 83298 115726 83310 115778
rect 110114 115726 110126 115778
rect 110178 115726 110190 115778
rect 111234 115726 111246 115778
rect 111298 115726 111310 115778
rect 117842 115726 117854 115778
rect 117906 115726 117918 115778
rect 10670 115714 10722 115726
rect 72606 115714 72658 115726
rect 10334 115666 10386 115678
rect 69022 115666 69074 115678
rect 3042 115614 3054 115666
rect 3106 115614 3118 115666
rect 4610 115614 4622 115666
rect 4674 115614 4686 115666
rect 11218 115614 11230 115666
rect 11282 115614 11294 115666
rect 23314 115614 23326 115666
rect 23378 115614 23390 115666
rect 32834 115614 32846 115666
rect 32898 115614 32910 115666
rect 36418 115614 36430 115666
rect 36482 115614 36494 115666
rect 47282 115614 47294 115666
rect 47346 115614 47358 115666
rect 56466 115614 56478 115666
rect 56530 115614 56542 115666
rect 57810 115614 57822 115666
rect 57874 115614 57886 115666
rect 59378 115614 59390 115666
rect 59442 115614 59454 115666
rect 63970 115614 63982 115666
rect 64034 115614 64046 115666
rect 66994 115614 67006 115666
rect 67058 115614 67070 115666
rect 10334 115602 10386 115614
rect 69022 115602 69074 115614
rect 71710 115666 71762 115678
rect 87950 115666 88002 115678
rect 72370 115614 72382 115666
rect 72434 115614 72446 115666
rect 73490 115614 73502 115666
rect 73554 115614 73566 115666
rect 76850 115614 76862 115666
rect 76914 115614 76926 115666
rect 80098 115614 80110 115666
rect 80162 115614 80174 115666
rect 86258 115614 86270 115666
rect 86322 115614 86334 115666
rect 101042 115614 101054 115666
rect 101106 115614 101118 115666
rect 112354 115614 112366 115666
rect 112418 115614 112430 115666
rect 116162 115614 116174 115666
rect 116226 115614 116238 115666
rect 116946 115614 116958 115666
rect 117010 115614 117022 115666
rect 71710 115602 71762 115614
rect 87950 115602 88002 115614
rect 5294 115554 5346 115566
rect 5294 115490 5346 115502
rect 9774 115554 9826 115566
rect 24670 115554 24722 115566
rect 33630 115554 33682 115566
rect 64430 115554 64482 115566
rect 11890 115502 11902 115554
rect 11954 115502 11966 115554
rect 14242 115502 14254 115554
rect 14306 115502 14318 115554
rect 30370 115502 30382 115554
rect 30434 115502 30446 115554
rect 32050 115502 32062 115554
rect 32114 115502 32126 115554
rect 38658 115502 38670 115554
rect 38722 115502 38734 115554
rect 44482 115502 44494 115554
rect 44546 115502 44558 115554
rect 46498 115502 46510 115554
rect 46562 115502 46574 115554
rect 47954 115502 47966 115554
rect 48018 115502 48030 115554
rect 55682 115502 55694 115554
rect 55746 115502 55758 115554
rect 58258 115502 58270 115554
rect 58322 115502 58334 115554
rect 60050 115502 60062 115554
rect 60114 115502 60126 115554
rect 9774 115490 9826 115502
rect 24670 115490 24722 115502
rect 33630 115490 33682 115502
rect 64430 115490 64482 115502
rect 66334 115554 66386 115566
rect 66334 115490 66386 115502
rect 70142 115554 70194 115566
rect 70142 115490 70194 115502
rect 71262 115554 71314 115566
rect 76414 115554 76466 115566
rect 80558 115554 80610 115566
rect 84142 115554 84194 115566
rect 74162 115502 74174 115554
rect 74226 115502 74238 115554
rect 77522 115502 77534 115554
rect 77586 115502 77598 115554
rect 82226 115502 82238 115554
rect 82290 115502 82302 115554
rect 71262 115490 71314 115502
rect 76414 115490 76466 115502
rect 80558 115490 80610 115502
rect 84142 115490 84194 115502
rect 85822 115554 85874 115566
rect 100494 115554 100546 115566
rect 86930 115502 86942 115554
rect 86994 115502 87006 115554
rect 101714 115502 101726 115554
rect 101778 115502 101790 115554
rect 109106 115502 109118 115554
rect 109170 115502 109182 115554
rect 115490 115502 115502 115554
rect 115554 115502 115566 115554
rect 85822 115490 85874 115502
rect 100494 115490 100546 115502
rect 1344 115274 118608 115308
rect 1344 115222 4478 115274
rect 4530 115222 4582 115274
rect 4634 115222 4686 115274
rect 4738 115222 35198 115274
rect 35250 115222 35302 115274
rect 35354 115222 35406 115274
rect 35458 115222 65918 115274
rect 65970 115222 66022 115274
rect 66074 115222 66126 115274
rect 66178 115222 96638 115274
rect 96690 115222 96742 115274
rect 96794 115222 96846 115274
rect 96898 115222 118608 115274
rect 1344 115188 118608 115222
rect 4398 114994 4450 115006
rect 2034 114942 2046 114994
rect 2098 114942 2110 114994
rect 4398 114930 4450 114942
rect 11342 114994 11394 115006
rect 11342 114930 11394 114942
rect 12350 114994 12402 115006
rect 36654 114994 36706 115006
rect 33954 114942 33966 114994
rect 34018 114942 34030 114994
rect 12350 114930 12402 114942
rect 36654 114930 36706 114942
rect 45390 114994 45442 115006
rect 45390 114930 45442 114942
rect 46958 114994 47010 115006
rect 46958 114930 47010 114942
rect 59166 114994 59218 115006
rect 59166 114930 59218 114942
rect 62974 114994 63026 115006
rect 62974 114930 63026 114942
rect 72158 114994 72210 115006
rect 72158 114930 72210 114942
rect 77870 114994 77922 115006
rect 115826 114942 115838 114994
rect 115890 114942 115902 114994
rect 77870 114930 77922 114942
rect 3614 114882 3666 114894
rect 3042 114830 3054 114882
rect 3106 114830 3118 114882
rect 3614 114818 3666 114830
rect 11902 114882 11954 114894
rect 64430 114882 64482 114894
rect 34850 114830 34862 114882
rect 34914 114830 34926 114882
rect 63634 114830 63646 114882
rect 63698 114830 63710 114882
rect 11902 114818 11954 114830
rect 64430 114818 64482 114830
rect 110798 114882 110850 114894
rect 110798 114818 110850 114830
rect 114382 114882 114434 114894
rect 115154 114830 115166 114882
rect 115218 114830 115230 114882
rect 117282 114830 117294 114882
rect 117346 114830 117358 114882
rect 114382 114818 114434 114830
rect 3950 114770 4002 114782
rect 3950 114706 4002 114718
rect 56926 114770 56978 114782
rect 56926 114706 56978 114718
rect 57486 114770 57538 114782
rect 57486 114706 57538 114718
rect 57822 114770 57874 114782
rect 57822 114706 57874 114718
rect 63870 114770 63922 114782
rect 86942 114770 86994 114782
rect 64754 114718 64766 114770
rect 64818 114718 64830 114770
rect 63870 114706 63922 114718
rect 86942 114706 86994 114718
rect 117070 114770 117122 114782
rect 117070 114706 117122 114718
rect 23774 114658 23826 114670
rect 23774 114594 23826 114606
rect 35534 114658 35586 114670
rect 35534 114594 35586 114606
rect 56478 114658 56530 114670
rect 56478 114594 56530 114606
rect 1344 114490 118608 114524
rect 1344 114438 19838 114490
rect 19890 114438 19942 114490
rect 19994 114438 20046 114490
rect 20098 114438 50558 114490
rect 50610 114438 50662 114490
rect 50714 114438 50766 114490
rect 50818 114438 81278 114490
rect 81330 114438 81382 114490
rect 81434 114438 81486 114490
rect 81538 114438 111998 114490
rect 112050 114438 112102 114490
rect 112154 114438 112206 114490
rect 112258 114438 118608 114490
rect 1344 114404 118608 114438
rect 64094 114322 64146 114334
rect 64094 114258 64146 114270
rect 117070 114322 117122 114334
rect 117070 114258 117122 114270
rect 1922 114158 1934 114210
rect 1986 114158 1998 114210
rect 3726 114098 3778 114110
rect 116162 114046 116174 114098
rect 116226 114046 116238 114098
rect 3726 114034 3778 114046
rect 116734 113986 116786 113998
rect 3266 113934 3278 113986
rect 3330 113934 3342 113986
rect 115490 113934 115502 113986
rect 115554 113934 115566 113986
rect 116162 113934 116174 113986
rect 116226 113983 116238 113986
rect 116226 113937 116447 113983
rect 116226 113934 116238 113937
rect 116401 113871 116447 113937
rect 116734 113922 116786 113934
rect 116722 113871 116734 113874
rect 116401 113825 116734 113871
rect 116722 113822 116734 113825
rect 116786 113822 116798 113874
rect 1344 113706 118608 113740
rect 1344 113654 4478 113706
rect 4530 113654 4582 113706
rect 4634 113654 4686 113706
rect 4738 113654 35198 113706
rect 35250 113654 35302 113706
rect 35354 113654 35406 113706
rect 35458 113654 65918 113706
rect 65970 113654 66022 113706
rect 66074 113654 66126 113706
rect 66178 113654 96638 113706
rect 96690 113654 96742 113706
rect 96794 113654 96846 113706
rect 96898 113654 118608 113706
rect 1344 113620 118608 113654
rect 1822 113426 1874 113438
rect 1822 113362 1874 113374
rect 2830 113202 2882 113214
rect 2830 113138 2882 113150
rect 2494 113090 2546 113102
rect 2494 113026 2546 113038
rect 3278 113090 3330 113102
rect 3278 113026 3330 113038
rect 1344 112922 118608 112956
rect 1344 112870 19838 112922
rect 19890 112870 19942 112922
rect 19994 112870 20046 112922
rect 20098 112870 50558 112922
rect 50610 112870 50662 112922
rect 50714 112870 50766 112922
rect 50818 112870 81278 112922
rect 81330 112870 81382 112922
rect 81434 112870 81486 112922
rect 81538 112870 111998 112922
rect 112050 112870 112102 112922
rect 112154 112870 112206 112922
rect 112258 112870 118608 112922
rect 1344 112836 118608 112870
rect 118078 112642 118130 112654
rect 118078 112578 118130 112590
rect 2818 112478 2830 112530
rect 2882 112478 2894 112530
rect 1922 112366 1934 112418
rect 1986 112366 1998 112418
rect 1344 112138 118608 112172
rect 1344 112086 4478 112138
rect 4530 112086 4582 112138
rect 4634 112086 4686 112138
rect 4738 112086 35198 112138
rect 35250 112086 35302 112138
rect 35354 112086 35406 112138
rect 35458 112086 65918 112138
rect 65970 112086 66022 112138
rect 66074 112086 66126 112138
rect 66178 112086 96638 112138
rect 96690 112086 96742 112138
rect 96794 112086 96846 112138
rect 96898 112086 118608 112138
rect 1344 112052 118608 112086
rect 3266 111806 3278 111858
rect 3330 111806 3342 111858
rect 1922 111582 1934 111634
rect 1986 111582 1998 111634
rect 118078 111522 118130 111534
rect 118078 111458 118130 111470
rect 1344 111354 118608 111388
rect 1344 111302 19838 111354
rect 19890 111302 19942 111354
rect 19994 111302 20046 111354
rect 20098 111302 50558 111354
rect 50610 111302 50662 111354
rect 50714 111302 50766 111354
rect 50818 111302 81278 111354
rect 81330 111302 81382 111354
rect 81434 111302 81486 111354
rect 81538 111302 111998 111354
rect 112050 111302 112102 111354
rect 112154 111302 112206 111354
rect 112258 111302 118608 111354
rect 1344 111268 118608 111302
rect 1710 111074 1762 111086
rect 1710 111010 1762 111022
rect 115154 110910 115166 110962
rect 115218 110910 115230 110962
rect 116622 110850 116674 110862
rect 115826 110798 115838 110850
rect 115890 110798 115902 110850
rect 116622 110786 116674 110798
rect 1344 110570 118608 110604
rect 1344 110518 4478 110570
rect 4530 110518 4582 110570
rect 4634 110518 4686 110570
rect 4738 110518 35198 110570
rect 35250 110518 35302 110570
rect 35354 110518 35406 110570
rect 35458 110518 65918 110570
rect 65970 110518 66022 110570
rect 66074 110518 66126 110570
rect 66178 110518 96638 110570
rect 96690 110518 96742 110570
rect 96794 110518 96846 110570
rect 96898 110518 118608 110570
rect 1344 110484 118608 110518
rect 1822 109954 1874 109966
rect 1822 109890 1874 109902
rect 1344 109786 118608 109820
rect 1344 109734 19838 109786
rect 19890 109734 19942 109786
rect 19994 109734 20046 109786
rect 20098 109734 50558 109786
rect 50610 109734 50662 109786
rect 50714 109734 50766 109786
rect 50818 109734 81278 109786
rect 81330 109734 81382 109786
rect 81434 109734 81486 109786
rect 81538 109734 111998 109786
rect 112050 109734 112102 109786
rect 112154 109734 112206 109786
rect 112258 109734 118608 109786
rect 1344 109700 118608 109734
rect 116274 109454 116286 109506
rect 116338 109454 116350 109506
rect 116846 109282 116898 109294
rect 114930 109230 114942 109282
rect 114994 109230 115006 109282
rect 116846 109218 116898 109230
rect 1344 109002 118608 109036
rect 1344 108950 4478 109002
rect 4530 108950 4582 109002
rect 4634 108950 4686 109002
rect 4738 108950 35198 109002
rect 35250 108950 35302 109002
rect 35354 108950 35406 109002
rect 35458 108950 65918 109002
rect 65970 108950 66022 109002
rect 66074 108950 66126 109002
rect 66178 108950 96638 109002
rect 96690 108950 96742 109002
rect 96794 108950 96846 109002
rect 96898 108950 118608 109002
rect 1344 108916 118608 108950
rect 1344 108218 118608 108252
rect 1344 108166 19838 108218
rect 19890 108166 19942 108218
rect 19994 108166 20046 108218
rect 20098 108166 50558 108218
rect 50610 108166 50662 108218
rect 50714 108166 50766 108218
rect 50818 108166 81278 108218
rect 81330 108166 81382 108218
rect 81434 108166 81486 108218
rect 81538 108166 111998 108218
rect 112050 108166 112102 108218
rect 112154 108166 112206 108218
rect 112258 108166 118608 108218
rect 1344 108132 118608 108166
rect 1822 107938 1874 107950
rect 116274 107886 116286 107938
rect 116338 107886 116350 107938
rect 1822 107874 1874 107886
rect 116846 107714 116898 107726
rect 114930 107662 114942 107714
rect 114994 107662 115006 107714
rect 116846 107650 116898 107662
rect 1344 107434 118608 107468
rect 1344 107382 4478 107434
rect 4530 107382 4582 107434
rect 4634 107382 4686 107434
rect 4738 107382 35198 107434
rect 35250 107382 35302 107434
rect 35354 107382 35406 107434
rect 35458 107382 65918 107434
rect 65970 107382 66022 107434
rect 66074 107382 66126 107434
rect 66178 107382 96638 107434
rect 96690 107382 96742 107434
rect 96794 107382 96846 107434
rect 96898 107382 118608 107434
rect 1344 107348 118608 107382
rect 118078 106818 118130 106830
rect 118078 106754 118130 106766
rect 1344 106650 118608 106684
rect 1344 106598 19838 106650
rect 19890 106598 19942 106650
rect 19994 106598 20046 106650
rect 20098 106598 50558 106650
rect 50610 106598 50662 106650
rect 50714 106598 50766 106650
rect 50818 106598 81278 106650
rect 81330 106598 81382 106650
rect 81434 106598 81486 106650
rect 81538 106598 111998 106650
rect 112050 106598 112102 106650
rect 112154 106598 112206 106650
rect 112258 106598 118608 106650
rect 1344 106564 118608 106598
rect 114494 106258 114546 106270
rect 114930 106206 114942 106258
rect 114994 106206 115006 106258
rect 114494 106194 114546 106206
rect 115826 106094 115838 106146
rect 115890 106094 115902 106146
rect 1344 105866 118608 105900
rect 1344 105814 4478 105866
rect 4530 105814 4582 105866
rect 4634 105814 4686 105866
rect 4738 105814 35198 105866
rect 35250 105814 35302 105866
rect 35354 105814 35406 105866
rect 35458 105814 65918 105866
rect 65970 105814 66022 105866
rect 66074 105814 66126 105866
rect 66178 105814 96638 105866
rect 96690 105814 96742 105866
rect 96794 105814 96846 105866
rect 96898 105814 118608 105866
rect 1344 105780 118608 105814
rect 1344 105082 118608 105116
rect 1344 105030 19838 105082
rect 19890 105030 19942 105082
rect 19994 105030 20046 105082
rect 20098 105030 50558 105082
rect 50610 105030 50662 105082
rect 50714 105030 50766 105082
rect 50818 105030 81278 105082
rect 81330 105030 81382 105082
rect 81434 105030 81486 105082
rect 81538 105030 111998 105082
rect 112050 105030 112102 105082
rect 112154 105030 112206 105082
rect 112258 105030 118608 105082
rect 1344 104996 118608 105030
rect 116274 104750 116286 104802
rect 116338 104750 116350 104802
rect 3042 104638 3054 104690
rect 3106 104638 3118 104690
rect 3614 104578 3666 104590
rect 116846 104578 116898 104590
rect 1922 104526 1934 104578
rect 1986 104526 1998 104578
rect 114930 104526 114942 104578
rect 114994 104526 115006 104578
rect 3614 104514 3666 104526
rect 116846 104514 116898 104526
rect 1344 104298 118608 104332
rect 1344 104246 4478 104298
rect 4530 104246 4582 104298
rect 4634 104246 4686 104298
rect 4738 104246 35198 104298
rect 35250 104246 35302 104298
rect 35354 104246 35406 104298
rect 35458 104246 65918 104298
rect 65970 104246 66022 104298
rect 66074 104246 66126 104298
rect 66178 104246 96638 104298
rect 96690 104246 96742 104298
rect 96794 104246 96846 104298
rect 96898 104246 118608 104298
rect 1344 104212 118608 104246
rect 1344 103514 118608 103548
rect 1344 103462 19838 103514
rect 19890 103462 19942 103514
rect 19994 103462 20046 103514
rect 20098 103462 50558 103514
rect 50610 103462 50662 103514
rect 50714 103462 50766 103514
rect 50818 103462 81278 103514
rect 81330 103462 81382 103514
rect 81434 103462 81486 103514
rect 81538 103462 111998 103514
rect 112050 103462 112102 103514
rect 112154 103462 112206 103514
rect 112258 103462 118608 103514
rect 1344 103428 118608 103462
rect 44830 103234 44882 103246
rect 44830 103170 44882 103182
rect 45166 103122 45218 103134
rect 3042 103070 3054 103122
rect 3106 103070 3118 103122
rect 45166 103058 45218 103070
rect 3614 103010 3666 103022
rect 1922 102958 1934 103010
rect 1986 102958 1998 103010
rect 3614 102946 3666 102958
rect 45614 103010 45666 103022
rect 45614 102946 45666 102958
rect 1344 102730 118608 102764
rect 1344 102678 4478 102730
rect 4530 102678 4582 102730
rect 4634 102678 4686 102730
rect 4738 102678 35198 102730
rect 35250 102678 35302 102730
rect 35354 102678 35406 102730
rect 35458 102678 65918 102730
rect 65970 102678 66022 102730
rect 66074 102678 66126 102730
rect 66178 102678 96638 102730
rect 96690 102678 96742 102730
rect 96794 102678 96846 102730
rect 96898 102678 118608 102730
rect 1344 102644 118608 102678
rect 3154 102398 3166 102450
rect 3218 102398 3230 102450
rect 114818 102398 114830 102450
rect 114882 102398 114894 102450
rect 2258 102174 2270 102226
rect 2322 102174 2334 102226
rect 116050 102174 116062 102226
rect 116114 102174 116126 102226
rect 117070 102114 117122 102126
rect 117070 102050 117122 102062
rect 1344 101946 118608 101980
rect 1344 101894 19838 101946
rect 19890 101894 19942 101946
rect 19994 101894 20046 101946
rect 20098 101894 50558 101946
rect 50610 101894 50662 101946
rect 50714 101894 50766 101946
rect 50818 101894 81278 101946
rect 81330 101894 81382 101946
rect 81434 101894 81486 101946
rect 81538 101894 111998 101946
rect 112050 101894 112102 101946
rect 112154 101894 112206 101946
rect 112258 101894 118608 101946
rect 1344 101860 118608 101894
rect 1822 101666 1874 101678
rect 1822 101602 1874 101614
rect 2382 101666 2434 101678
rect 2382 101602 2434 101614
rect 118078 101666 118130 101678
rect 118078 101602 118130 101614
rect 1344 101162 118608 101196
rect 1344 101110 4478 101162
rect 4530 101110 4582 101162
rect 4634 101110 4686 101162
rect 4738 101110 35198 101162
rect 35250 101110 35302 101162
rect 35354 101110 35406 101162
rect 35458 101110 65918 101162
rect 65970 101110 66022 101162
rect 66074 101110 66126 101162
rect 66178 101110 96638 101162
rect 96690 101110 96742 101162
rect 96794 101110 96846 101162
rect 96898 101110 118608 101162
rect 1344 101076 118608 101110
rect 1344 100378 118608 100412
rect 1344 100326 19838 100378
rect 19890 100326 19942 100378
rect 19994 100326 20046 100378
rect 20098 100326 50558 100378
rect 50610 100326 50662 100378
rect 50714 100326 50766 100378
rect 50818 100326 81278 100378
rect 81330 100326 81382 100378
rect 81434 100326 81486 100378
rect 81538 100326 111998 100378
rect 112050 100326 112102 100378
rect 112154 100326 112206 100378
rect 112258 100326 118608 100378
rect 1344 100292 118608 100326
rect 1922 100046 1934 100098
rect 1986 100046 1998 100098
rect 114494 99986 114546 99998
rect 114930 99934 114942 99986
rect 114994 99934 115006 99986
rect 114494 99922 114546 99934
rect 3266 99822 3278 99874
rect 3330 99822 3342 99874
rect 115826 99822 115838 99874
rect 115890 99822 115902 99874
rect 1344 99594 118608 99628
rect 1344 99542 4478 99594
rect 4530 99542 4582 99594
rect 4634 99542 4686 99594
rect 4738 99542 35198 99594
rect 35250 99542 35302 99594
rect 35354 99542 35406 99594
rect 35458 99542 65918 99594
rect 65970 99542 66022 99594
rect 66074 99542 66126 99594
rect 66178 99542 96638 99594
rect 96690 99542 96742 99594
rect 96794 99542 96846 99594
rect 96898 99542 118608 99594
rect 1344 99508 118608 99542
rect 38558 99426 38610 99438
rect 38558 99362 38610 99374
rect 1822 99314 1874 99326
rect 1822 99250 1874 99262
rect 37886 99314 37938 99326
rect 37886 99250 37938 99262
rect 38334 99314 38386 99326
rect 38334 99250 38386 99262
rect 39454 99314 39506 99326
rect 39454 99250 39506 99262
rect 2594 99150 2606 99202
rect 2658 99150 2670 99202
rect 38882 99150 38894 99202
rect 38946 99150 38958 99202
rect 2830 98978 2882 98990
rect 2830 98914 2882 98926
rect 3278 98978 3330 98990
rect 3278 98914 3330 98926
rect 1344 98810 118608 98844
rect 1344 98758 19838 98810
rect 19890 98758 19942 98810
rect 19994 98758 20046 98810
rect 20098 98758 50558 98810
rect 50610 98758 50662 98810
rect 50714 98758 50766 98810
rect 50818 98758 81278 98810
rect 81330 98758 81382 98810
rect 81434 98758 81486 98810
rect 81538 98758 111998 98810
rect 112050 98758 112102 98810
rect 112154 98758 112206 98810
rect 112258 98758 118608 98810
rect 1344 98724 118608 98758
rect 2818 98366 2830 98418
rect 2882 98366 2894 98418
rect 1922 98254 1934 98306
rect 1986 98254 1998 98306
rect 1344 98026 118608 98060
rect 1344 97974 4478 98026
rect 4530 97974 4582 98026
rect 4634 97974 4686 98026
rect 4738 97974 35198 98026
rect 35250 97974 35302 98026
rect 35354 97974 35406 98026
rect 35458 97974 65918 98026
rect 65970 97974 66022 98026
rect 66074 97974 66126 98026
rect 66178 97974 96638 98026
rect 96690 97974 96742 98026
rect 96794 97974 96846 98026
rect 96898 97974 118608 98026
rect 1344 97940 118608 97974
rect 3266 97694 3278 97746
rect 3330 97694 3342 97746
rect 1922 97470 1934 97522
rect 1986 97470 1998 97522
rect 1344 97242 118608 97276
rect 1344 97190 19838 97242
rect 19890 97190 19942 97242
rect 19994 97190 20046 97242
rect 20098 97190 50558 97242
rect 50610 97190 50662 97242
rect 50714 97190 50766 97242
rect 50818 97190 81278 97242
rect 81330 97190 81382 97242
rect 81434 97190 81486 97242
rect 81538 97190 111998 97242
rect 112050 97190 112102 97242
rect 112154 97190 112206 97242
rect 112258 97190 118608 97242
rect 1344 97156 118608 97190
rect 1710 96962 1762 96974
rect 1710 96898 1762 96910
rect 118078 96962 118130 96974
rect 118078 96898 118130 96910
rect 1344 96458 118608 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 65918 96458
rect 65970 96406 66022 96458
rect 66074 96406 66126 96458
rect 66178 96406 96638 96458
rect 96690 96406 96742 96458
rect 96794 96406 96846 96458
rect 96898 96406 118608 96458
rect 1344 96372 118608 96406
rect 1344 95674 118608 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 50558 95674
rect 50610 95622 50662 95674
rect 50714 95622 50766 95674
rect 50818 95622 81278 95674
rect 81330 95622 81382 95674
rect 81434 95622 81486 95674
rect 81538 95622 111998 95674
rect 112050 95622 112102 95674
rect 112154 95622 112206 95674
rect 112258 95622 118608 95674
rect 1344 95588 118608 95622
rect 2818 95230 2830 95282
rect 2882 95230 2894 95282
rect 114930 95230 114942 95282
rect 114994 95230 115006 95282
rect 114494 95170 114546 95182
rect 1922 95118 1934 95170
rect 1986 95118 1998 95170
rect 115826 95118 115838 95170
rect 115890 95118 115902 95170
rect 114494 95106 114546 95118
rect 1344 94890 118608 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 65918 94890
rect 65970 94838 66022 94890
rect 66074 94838 66126 94890
rect 66178 94838 96638 94890
rect 96690 94838 96742 94890
rect 96794 94838 96846 94890
rect 96898 94838 118608 94890
rect 1344 94804 118608 94838
rect 3278 94610 3330 94622
rect 114818 94558 114830 94610
rect 114882 94558 114894 94610
rect 3278 94546 3330 94558
rect 2830 94498 2882 94510
rect 2830 94434 2882 94446
rect 2494 94386 2546 94398
rect 2494 94322 2546 94334
rect 71262 94386 71314 94398
rect 71262 94322 71314 94334
rect 71822 94386 71874 94398
rect 116050 94334 116062 94386
rect 116114 94334 116126 94386
rect 71822 94322 71874 94334
rect 72158 94274 72210 94286
rect 72158 94210 72210 94222
rect 117070 94274 117122 94286
rect 117070 94210 117122 94222
rect 1344 94106 118608 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 50558 94106
rect 50610 94054 50662 94106
rect 50714 94054 50766 94106
rect 50818 94054 81278 94106
rect 81330 94054 81382 94106
rect 81434 94054 81486 94106
rect 81538 94054 111998 94106
rect 112050 94054 112102 94106
rect 112154 94054 112206 94106
rect 112258 94054 118608 94106
rect 1344 94020 118608 94054
rect 48302 93826 48354 93838
rect 48302 93762 48354 93774
rect 48638 93714 48690 93726
rect 3042 93662 3054 93714
rect 3106 93662 3118 93714
rect 48638 93650 48690 93662
rect 3614 93602 3666 93614
rect 1922 93550 1934 93602
rect 1986 93550 1998 93602
rect 3614 93538 3666 93550
rect 49422 93602 49474 93614
rect 49422 93538 49474 93550
rect 1344 93322 118608 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 65918 93322
rect 65970 93270 66022 93322
rect 66074 93270 66126 93322
rect 66178 93270 96638 93322
rect 96690 93270 96742 93322
rect 96794 93270 96846 93322
rect 96898 93270 118608 93322
rect 1344 93236 118608 93270
rect 3266 92990 3278 93042
rect 3330 92990 3342 93042
rect 115826 92990 115838 93042
rect 115890 92990 115902 93042
rect 114382 92930 114434 92942
rect 114930 92878 114942 92930
rect 114994 92878 115006 92930
rect 114382 92866 114434 92878
rect 1922 92766 1934 92818
rect 1986 92766 1998 92818
rect 1344 92538 118608 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 50558 92538
rect 50610 92486 50662 92538
rect 50714 92486 50766 92538
rect 50818 92486 81278 92538
rect 81330 92486 81382 92538
rect 81434 92486 81486 92538
rect 81538 92486 111998 92538
rect 112050 92486 112102 92538
rect 112154 92486 112206 92538
rect 112258 92486 118608 92538
rect 1344 92452 118608 92486
rect 1822 92370 1874 92382
rect 1822 92306 1874 92318
rect 1344 91754 118608 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 65918 91754
rect 65970 91702 66022 91754
rect 66074 91702 66126 91754
rect 66178 91702 96638 91754
rect 96690 91702 96742 91754
rect 96794 91702 96846 91754
rect 96898 91702 118608 91754
rect 1344 91668 118608 91702
rect 1344 90970 118608 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 50558 90970
rect 50610 90918 50662 90970
rect 50714 90918 50766 90970
rect 50818 90918 81278 90970
rect 81330 90918 81382 90970
rect 81434 90918 81486 90970
rect 81538 90918 111998 90970
rect 112050 90918 112102 90970
rect 112154 90918 112206 90970
rect 112258 90918 118608 90970
rect 1344 90884 118608 90918
rect 2818 90526 2830 90578
rect 2882 90526 2894 90578
rect 1922 90414 1934 90466
rect 1986 90414 1998 90466
rect 1344 90186 118608 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 65918 90186
rect 65970 90134 66022 90186
rect 66074 90134 66126 90186
rect 66178 90134 96638 90186
rect 96690 90134 96742 90186
rect 96794 90134 96846 90186
rect 96898 90134 118608 90186
rect 1344 90100 118608 90134
rect 3042 89966 3054 90018
rect 3106 90015 3118 90018
rect 3266 90015 3278 90018
rect 3106 89969 3278 90015
rect 3106 89966 3118 89969
rect 3266 89966 3278 89969
rect 3330 89966 3342 90018
rect 3278 89906 3330 89918
rect 115378 89854 115390 89906
rect 115442 89854 115454 89906
rect 3278 89842 3330 89854
rect 2830 89794 2882 89806
rect 115938 89742 115950 89794
rect 116002 89742 116014 89794
rect 2830 89730 2882 89742
rect 2494 89682 2546 89694
rect 2494 89618 2546 89630
rect 58830 89682 58882 89694
rect 58830 89618 58882 89630
rect 59166 89682 59218 89694
rect 59166 89618 59218 89630
rect 116958 89682 117010 89694
rect 116958 89618 117010 89630
rect 59726 89570 59778 89582
rect 59726 89506 59778 89518
rect 1344 89402 118608 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 50558 89402
rect 50610 89350 50662 89402
rect 50714 89350 50766 89402
rect 50818 89350 81278 89402
rect 81330 89350 81382 89402
rect 81434 89350 81486 89402
rect 81538 89350 111998 89402
rect 112050 89350 112102 89402
rect 112154 89350 112206 89402
rect 112258 89350 118608 89402
rect 1344 89316 118608 89350
rect 3502 89010 3554 89022
rect 3042 88958 3054 89010
rect 3106 88958 3118 89010
rect 3502 88946 3554 88958
rect 1922 88846 1934 88898
rect 1986 88846 1998 88898
rect 1344 88618 118608 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 65918 88618
rect 65970 88566 66022 88618
rect 66074 88566 66126 88618
rect 66178 88566 96638 88618
rect 96690 88566 96742 88618
rect 96794 88566 96846 88618
rect 96898 88566 118608 88618
rect 1344 88532 118608 88566
rect 3266 88286 3278 88338
rect 3330 88286 3342 88338
rect 1922 88062 1934 88114
rect 1986 88062 1998 88114
rect 1344 87834 118608 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 50558 87834
rect 50610 87782 50662 87834
rect 50714 87782 50766 87834
rect 50818 87782 81278 87834
rect 81330 87782 81382 87834
rect 81434 87782 81486 87834
rect 81538 87782 111998 87834
rect 112050 87782 112102 87834
rect 112154 87782 112206 87834
rect 112258 87782 118608 87834
rect 1344 87748 118608 87782
rect 1822 87666 1874 87678
rect 1822 87602 1874 87614
rect 116274 87502 116286 87554
rect 116338 87502 116350 87554
rect 116846 87442 116898 87454
rect 116846 87378 116898 87390
rect 114930 87278 114942 87330
rect 114994 87278 115006 87330
rect 1344 87050 118608 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 65918 87050
rect 65970 86998 66022 87050
rect 66074 86998 66126 87050
rect 66178 86998 96638 87050
rect 96690 86998 96742 87050
rect 96794 86998 96846 87050
rect 96898 86998 118608 87050
rect 1344 86964 118608 86998
rect 115826 86718 115838 86770
rect 115890 86718 115902 86770
rect 114382 86658 114434 86670
rect 114930 86606 114942 86658
rect 114994 86606 115006 86658
rect 114382 86594 114434 86606
rect 1344 86266 118608 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 50558 86266
rect 50610 86214 50662 86266
rect 50714 86214 50766 86266
rect 50818 86214 81278 86266
rect 81330 86214 81382 86266
rect 81434 86214 81486 86266
rect 81538 86214 111998 86266
rect 112050 86214 112102 86266
rect 112154 86214 112206 86266
rect 112258 86214 118608 86266
rect 1344 86180 118608 86214
rect 1822 85986 1874 85998
rect 1822 85922 1874 85934
rect 1344 85482 118608 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 65918 85482
rect 65970 85430 66022 85482
rect 66074 85430 66126 85482
rect 66178 85430 96638 85482
rect 96690 85430 96742 85482
rect 96794 85430 96846 85482
rect 96898 85430 118608 85482
rect 1344 85396 118608 85430
rect 115826 85150 115838 85202
rect 115890 85150 115902 85202
rect 114494 85090 114546 85102
rect 114930 85038 114942 85090
rect 114994 85038 115006 85090
rect 114494 85026 114546 85038
rect 76190 84978 76242 84990
rect 76190 84914 76242 84926
rect 75630 84866 75682 84878
rect 75630 84802 75682 84814
rect 76526 84866 76578 84878
rect 76526 84802 76578 84814
rect 1344 84698 118608 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 50558 84698
rect 50610 84646 50662 84698
rect 50714 84646 50766 84698
rect 50818 84646 81278 84698
rect 81330 84646 81382 84698
rect 81434 84646 81486 84698
rect 81538 84646 111998 84698
rect 112050 84646 112102 84698
rect 112154 84646 112206 84698
rect 112258 84646 118608 84698
rect 1344 84612 118608 84646
rect 1822 84418 1874 84430
rect 1822 84354 1874 84366
rect 1344 83914 118608 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 65918 83914
rect 65970 83862 66022 83914
rect 66074 83862 66126 83914
rect 66178 83862 96638 83914
rect 96690 83862 96742 83914
rect 96794 83862 96846 83914
rect 96898 83862 118608 83914
rect 1344 83828 118608 83862
rect 115378 83582 115390 83634
rect 115442 83582 115454 83634
rect 116162 83470 116174 83522
rect 116226 83470 116238 83522
rect 117282 83470 117294 83522
rect 117346 83470 117358 83522
rect 117070 83410 117122 83422
rect 117070 83346 117122 83358
rect 1344 83130 118608 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 50558 83130
rect 50610 83078 50662 83130
rect 50714 83078 50766 83130
rect 50818 83078 81278 83130
rect 81330 83078 81382 83130
rect 81434 83078 81486 83130
rect 81538 83078 111998 83130
rect 112050 83078 112102 83130
rect 112154 83078 112206 83130
rect 112258 83078 118608 83130
rect 1344 83044 118608 83078
rect 116734 82962 116786 82974
rect 116734 82898 116786 82910
rect 118078 82850 118130 82862
rect 118078 82786 118130 82798
rect 2818 82686 2830 82738
rect 2882 82686 2894 82738
rect 1922 82574 1934 82626
rect 1986 82574 1998 82626
rect 1344 82346 118608 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 65918 82346
rect 65970 82294 66022 82346
rect 66074 82294 66126 82346
rect 66178 82294 96638 82346
rect 96690 82294 96742 82346
rect 96794 82294 96846 82346
rect 96898 82294 118608 82346
rect 1344 82260 118608 82294
rect 3042 82126 3054 82178
rect 3106 82175 3118 82178
rect 3266 82175 3278 82178
rect 3106 82129 3278 82175
rect 3106 82126 3118 82129
rect 3266 82126 3278 82129
rect 3330 82126 3342 82178
rect 3278 82066 3330 82078
rect 3278 82002 3330 82014
rect 2830 81954 2882 81966
rect 2830 81890 2882 81902
rect 2494 81842 2546 81854
rect 2494 81778 2546 81790
rect 1344 81562 118608 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 50558 81562
rect 50610 81510 50662 81562
rect 50714 81510 50766 81562
rect 50818 81510 81278 81562
rect 81330 81510 81382 81562
rect 81434 81510 81486 81562
rect 81538 81510 111998 81562
rect 112050 81510 112102 81562
rect 112154 81510 112206 81562
rect 112258 81510 118608 81562
rect 1344 81476 118608 81510
rect 1344 80778 118608 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 65918 80778
rect 65970 80726 66022 80778
rect 66074 80726 66126 80778
rect 66178 80726 96638 80778
rect 96690 80726 96742 80778
rect 96794 80726 96846 80778
rect 96898 80726 118608 80778
rect 1344 80692 118608 80726
rect 2818 80334 2830 80386
rect 2882 80334 2894 80386
rect 1922 80222 1934 80274
rect 1986 80222 1998 80274
rect 1344 79994 118608 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 50558 79994
rect 50610 79942 50662 79994
rect 50714 79942 50766 79994
rect 50818 79942 81278 79994
rect 81330 79942 81382 79994
rect 81434 79942 81486 79994
rect 81538 79942 111998 79994
rect 112050 79942 112102 79994
rect 112154 79942 112206 79994
rect 112258 79942 118608 79994
rect 1344 79908 118608 79942
rect 2494 79826 2546 79838
rect 2494 79762 2546 79774
rect 3278 79826 3330 79838
rect 3278 79762 3330 79774
rect 117966 79826 118018 79838
rect 117966 79762 118018 79774
rect 117282 79662 117294 79714
rect 117346 79662 117358 79714
rect 2830 79602 2882 79614
rect 2830 79538 2882 79550
rect 114830 79378 114882 79390
rect 3042 79326 3054 79378
rect 3106 79375 3118 79378
rect 3266 79375 3278 79378
rect 3106 79329 3278 79375
rect 3106 79326 3118 79329
rect 3266 79326 3278 79329
rect 3330 79326 3342 79378
rect 114830 79314 114882 79326
rect 1344 79210 118608 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 65918 79210
rect 65970 79158 66022 79210
rect 66074 79158 66126 79210
rect 66178 79158 96638 79210
rect 96690 79158 96742 79210
rect 96794 79158 96846 79210
rect 96898 79158 118608 79210
rect 1344 79124 118608 79158
rect 3042 78766 3054 78818
rect 3106 78766 3118 78818
rect 1922 78654 1934 78706
rect 1986 78654 1998 78706
rect 3502 78594 3554 78606
rect 3502 78530 3554 78542
rect 118078 78594 118130 78606
rect 118078 78530 118130 78542
rect 1344 78426 118608 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 50558 78426
rect 50610 78374 50662 78426
rect 50714 78374 50766 78426
rect 50818 78374 81278 78426
rect 81330 78374 81382 78426
rect 81434 78374 81486 78426
rect 81538 78374 111998 78426
rect 112050 78374 112102 78426
rect 112154 78374 112206 78426
rect 112258 78374 118608 78426
rect 1344 78340 118608 78374
rect 117966 78258 118018 78270
rect 117966 78194 118018 78206
rect 117170 78094 117182 78146
rect 117234 78094 117246 78146
rect 114830 77810 114882 77822
rect 114830 77746 114882 77758
rect 1344 77642 118608 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 65918 77642
rect 65970 77590 66022 77642
rect 66074 77590 66126 77642
rect 66178 77590 96638 77642
rect 96690 77590 96742 77642
rect 96794 77590 96846 77642
rect 96898 77590 118608 77642
rect 1344 77556 118608 77590
rect 1822 77026 1874 77038
rect 1822 76962 1874 76974
rect 1344 76858 118608 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 81278 76858
rect 81330 76806 81382 76858
rect 81434 76806 81486 76858
rect 81538 76806 111998 76858
rect 112050 76806 112102 76858
rect 112154 76806 112206 76858
rect 112258 76806 118608 76858
rect 1344 76772 118608 76806
rect 1922 76526 1934 76578
rect 1986 76526 1998 76578
rect 4398 76242 4450 76254
rect 4398 76178 4450 76190
rect 1344 76074 118608 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 96638 76074
rect 96690 76022 96742 76074
rect 96794 76022 96846 76074
rect 96898 76022 118608 76074
rect 1344 75988 118608 76022
rect 114382 75682 114434 75694
rect 2818 75630 2830 75682
rect 2882 75630 2894 75682
rect 114930 75630 114942 75682
rect 114994 75630 115006 75682
rect 114382 75618 114434 75630
rect 1922 75518 1934 75570
rect 1986 75518 1998 75570
rect 116050 75518 116062 75570
rect 116114 75518 116126 75570
rect 1344 75290 118608 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 81278 75290
rect 81330 75238 81382 75290
rect 81434 75238 81486 75290
rect 81538 75238 111998 75290
rect 112050 75238 112102 75290
rect 112154 75238 112206 75290
rect 112258 75238 118608 75290
rect 1344 75204 118608 75238
rect 2494 75122 2546 75134
rect 2494 75058 2546 75070
rect 3278 75122 3330 75134
rect 3278 75058 3330 75070
rect 2830 75010 2882 75022
rect 2830 74946 2882 74958
rect 1344 74506 118608 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 96638 74506
rect 96690 74454 96742 74506
rect 96794 74454 96846 74506
rect 96898 74454 118608 74506
rect 1344 74420 118608 74454
rect 114818 74174 114830 74226
rect 114882 74174 114894 74226
rect 117070 74002 117122 74014
rect 116162 73950 116174 74002
rect 116226 73950 116238 74002
rect 117070 73938 117122 73950
rect 1344 73722 118608 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 81278 73722
rect 81330 73670 81382 73722
rect 81434 73670 81486 73722
rect 81538 73670 111998 73722
rect 112050 73670 112102 73722
rect 112154 73670 112206 73722
rect 112258 73670 118608 73722
rect 1344 73636 118608 73670
rect 1344 72938 118608 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 96638 72938
rect 96690 72886 96742 72938
rect 96794 72886 96846 72938
rect 96898 72886 118608 72938
rect 1344 72852 118608 72886
rect 1344 72154 118608 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 81278 72154
rect 81330 72102 81382 72154
rect 81434 72102 81486 72154
rect 81538 72102 111998 72154
rect 112050 72102 112102 72154
rect 112154 72102 112206 72154
rect 112258 72102 118608 72154
rect 1344 72068 118608 72102
rect 1922 71822 1934 71874
rect 1986 71822 1998 71874
rect 3266 71598 3278 71650
rect 3330 71598 3342 71650
rect 1344 71370 118608 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 96638 71370
rect 96690 71318 96742 71370
rect 96794 71318 96846 71370
rect 96898 71318 118608 71370
rect 1344 71284 118608 71318
rect 1822 71090 1874 71102
rect 1822 71026 1874 71038
rect 118078 70754 118130 70766
rect 118078 70690 118130 70702
rect 1344 70586 118608 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 81278 70586
rect 81330 70534 81382 70586
rect 81434 70534 81486 70586
rect 81538 70534 111998 70586
rect 112050 70534 112102 70586
rect 112154 70534 112206 70586
rect 112258 70534 118608 70586
rect 1344 70500 118608 70534
rect 3390 70418 3442 70430
rect 3390 70354 3442 70366
rect 115502 70418 115554 70430
rect 115502 70354 115554 70366
rect 115950 70418 116002 70430
rect 115950 70354 116002 70366
rect 2494 70306 2546 70318
rect 2494 70242 2546 70254
rect 2830 70306 2882 70318
rect 2830 70242 2882 70254
rect 1344 69802 118608 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 96638 69802
rect 96690 69750 96742 69802
rect 96794 69750 96846 69802
rect 96898 69750 118608 69802
rect 1344 69716 118608 69750
rect 115826 69470 115838 69522
rect 115890 69470 115902 69522
rect 114382 69410 114434 69422
rect 2818 69358 2830 69410
rect 2882 69358 2894 69410
rect 114930 69358 114942 69410
rect 114994 69358 115006 69410
rect 114382 69346 114434 69358
rect 1922 69246 1934 69298
rect 1986 69246 1998 69298
rect 55918 69186 55970 69198
rect 55918 69122 55970 69134
rect 117070 69186 117122 69198
rect 117070 69122 117122 69134
rect 1344 69018 118608 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 81278 69018
rect 81330 68966 81382 69018
rect 81434 68966 81486 69018
rect 81538 68966 111998 69018
rect 112050 68966 112102 69018
rect 112154 68966 112206 69018
rect 112258 68966 118608 69018
rect 1344 68932 118608 68966
rect 46398 68850 46450 68862
rect 46398 68786 46450 68798
rect 116386 68686 116398 68738
rect 116450 68686 116462 68738
rect 116946 68686 116958 68738
rect 117010 68686 117022 68738
rect 46062 68626 46114 68638
rect 3042 68574 3054 68626
rect 3106 68574 3118 68626
rect 114482 68574 114494 68626
rect 114546 68574 114558 68626
rect 46062 68562 46114 68574
rect 3614 68514 3666 68526
rect 1922 68462 1934 68514
rect 1986 68462 1998 68514
rect 3614 68450 3666 68462
rect 46846 68514 46898 68526
rect 46846 68450 46898 68462
rect 55246 68514 55298 68526
rect 55246 68450 55298 68462
rect 55694 68514 55746 68526
rect 55694 68450 55746 68462
rect 56142 68514 56194 68526
rect 56142 68450 56194 68462
rect 56478 68514 56530 68526
rect 56478 68450 56530 68462
rect 63086 68514 63138 68526
rect 63086 68450 63138 68462
rect 63982 68514 64034 68526
rect 63982 68450 64034 68462
rect 114046 68514 114098 68526
rect 115602 68462 115614 68514
rect 115666 68462 115678 68514
rect 114046 68450 114098 68462
rect 117182 68402 117234 68414
rect 117182 68338 117234 68350
rect 117518 68402 117570 68414
rect 117518 68338 117570 68350
rect 1344 68234 118608 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 96638 68234
rect 96690 68182 96742 68234
rect 96794 68182 96846 68234
rect 96898 68182 118608 68234
rect 1344 68148 118608 68182
rect 57026 68014 57038 68066
rect 57090 68014 57102 68066
rect 60622 67954 60674 67966
rect 64094 67954 64146 67966
rect 54898 67902 54910 67954
rect 54962 67902 54974 67954
rect 56578 67902 56590 67954
rect 56642 67902 56654 67954
rect 63634 67902 63646 67954
rect 63698 67902 63710 67954
rect 115490 67902 115502 67954
rect 115554 67902 115566 67954
rect 60622 67890 60674 67902
rect 64094 67890 64146 67902
rect 49310 67842 49362 67854
rect 61854 67842 61906 67854
rect 117406 67842 117458 67854
rect 55122 67790 55134 67842
rect 55186 67790 55198 67842
rect 56690 67790 56702 67842
rect 56754 67790 56766 67842
rect 62626 67790 62638 67842
rect 62690 67790 62702 67842
rect 74834 67790 74846 67842
rect 74898 67790 74910 67842
rect 77522 67790 77534 67842
rect 77586 67790 77598 67842
rect 116162 67790 116174 67842
rect 116226 67790 116238 67842
rect 49310 67778 49362 67790
rect 61854 67778 61906 67790
rect 117406 67778 117458 67790
rect 55694 67730 55746 67742
rect 63310 67730 63362 67742
rect 62514 67678 62526 67730
rect 62578 67678 62590 67730
rect 55694 67666 55746 67678
rect 63310 67666 63362 67678
rect 71710 67730 71762 67742
rect 71710 67666 71762 67678
rect 77758 67730 77810 67742
rect 77758 67666 77810 67678
rect 49646 67618 49698 67630
rect 49646 67554 49698 67566
rect 57822 67618 57874 67630
rect 57822 67554 57874 67566
rect 61518 67618 61570 67630
rect 61518 67554 61570 67566
rect 63534 67618 63586 67630
rect 63534 67554 63586 67566
rect 64542 67618 64594 67630
rect 64542 67554 64594 67566
rect 72046 67618 72098 67630
rect 72046 67554 72098 67566
rect 75070 67618 75122 67630
rect 75070 67554 75122 67566
rect 78318 67618 78370 67630
rect 78318 67554 78370 67566
rect 117070 67618 117122 67630
rect 117070 67554 117122 67566
rect 1344 67450 118608 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 81278 67450
rect 81330 67398 81382 67450
rect 81434 67398 81486 67450
rect 81538 67398 111998 67450
rect 112050 67398 112102 67450
rect 112154 67398 112206 67450
rect 112258 67398 118608 67450
rect 1344 67364 118608 67398
rect 56590 67282 56642 67294
rect 56590 67218 56642 67230
rect 71374 67282 71426 67294
rect 71374 67218 71426 67230
rect 82350 67282 82402 67294
rect 82350 67218 82402 67230
rect 48638 67170 48690 67182
rect 56254 67170 56306 67182
rect 50530 67118 50542 67170
rect 50594 67118 50606 67170
rect 48638 67106 48690 67118
rect 56254 67106 56306 67118
rect 56366 67170 56418 67182
rect 72258 67118 72270 67170
rect 72322 67118 72334 67170
rect 74946 67118 74958 67170
rect 75010 67118 75022 67170
rect 78418 67118 78430 67170
rect 78482 67118 78494 67170
rect 117282 67118 117294 67170
rect 117346 67118 117358 67170
rect 56366 67106 56418 67118
rect 49646 67058 49698 67070
rect 65326 67058 65378 67070
rect 82014 67058 82066 67070
rect 48402 67006 48414 67058
rect 48466 67006 48478 67058
rect 50754 67006 50766 67058
rect 50818 67006 50830 67058
rect 52658 67006 52670 67058
rect 52722 67006 52734 67058
rect 57586 67006 57598 67058
rect 57650 67006 57662 67058
rect 61282 67006 61294 67058
rect 61346 67006 61358 67058
rect 72370 67006 72382 67058
rect 72434 67006 72446 67058
rect 74274 67006 74286 67058
rect 74338 67006 74350 67058
rect 77634 67006 77646 67058
rect 77698 67006 77710 67058
rect 117954 67006 117966 67058
rect 118018 67006 118030 67058
rect 49646 66994 49698 67006
rect 65326 66994 65378 67006
rect 82014 66994 82066 67006
rect 51326 66946 51378 66958
rect 64542 66946 64594 66958
rect 53330 66894 53342 66946
rect 53394 66894 53406 66946
rect 55570 66894 55582 66946
rect 55634 66894 55646 66946
rect 58258 66894 58270 66946
rect 58322 66894 58334 66946
rect 60498 66894 60510 66946
rect 60562 66894 60574 66946
rect 61954 66894 61966 66946
rect 62018 66894 62030 66946
rect 64082 66894 64094 66946
rect 64146 66894 64158 66946
rect 51326 66882 51378 66894
rect 64542 66882 64594 66894
rect 70254 66946 70306 66958
rect 70254 66882 70306 66894
rect 70702 66946 70754 66958
rect 70702 66882 70754 66894
rect 73278 66946 73330 66958
rect 81230 66946 81282 66958
rect 77074 66894 77086 66946
rect 77138 66894 77150 66946
rect 80546 66894 80558 66946
rect 80610 66894 80622 66946
rect 73278 66882 73330 66894
rect 81230 66882 81282 66894
rect 113934 66946 113986 66958
rect 113934 66882 113986 66894
rect 114382 66946 114434 66958
rect 115154 66894 115166 66946
rect 115218 66894 115230 66946
rect 114382 66882 114434 66894
rect 49982 66834 50034 66846
rect 49982 66770 50034 66782
rect 71710 66834 71762 66846
rect 71710 66770 71762 66782
rect 1344 66666 118608 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 96638 66666
rect 96690 66614 96742 66666
rect 96794 66614 96846 66666
rect 96898 66614 118608 66666
rect 1344 66580 118608 66614
rect 53678 66498 53730 66510
rect 53678 66434 53730 66446
rect 74846 66498 74898 66510
rect 77870 66498 77922 66510
rect 76290 66446 76302 66498
rect 76354 66495 76366 66498
rect 76514 66495 76526 66498
rect 76354 66449 76526 66495
rect 76354 66446 76366 66449
rect 76514 66446 76526 66449
rect 76578 66446 76590 66498
rect 74846 66434 74898 66446
rect 77870 66434 77922 66446
rect 55470 66386 55522 66398
rect 3266 66334 3278 66386
rect 3330 66334 3342 66386
rect 47282 66334 47294 66386
rect 47346 66334 47358 66386
rect 49410 66334 49422 66386
rect 49474 66334 49486 66386
rect 55470 66322 55522 66334
rect 55918 66386 55970 66398
rect 55918 66322 55970 66334
rect 57262 66386 57314 66398
rect 57262 66322 57314 66334
rect 58270 66386 58322 66398
rect 58270 66322 58322 66334
rect 58942 66386 58994 66398
rect 58942 66322 58994 66334
rect 59390 66386 59442 66398
rect 59390 66322 59442 66334
rect 60622 66386 60674 66398
rect 76526 66386 76578 66398
rect 63746 66334 63758 66386
rect 63810 66334 63822 66386
rect 65874 66334 65886 66386
rect 65938 66334 65950 66386
rect 72034 66334 72046 66386
rect 72098 66334 72110 66386
rect 74162 66334 74174 66386
rect 74226 66334 74238 66386
rect 60622 66322 60674 66334
rect 76526 66322 76578 66334
rect 79550 66386 79602 66398
rect 79550 66322 79602 66334
rect 54798 66274 54850 66286
rect 45602 66222 45614 66274
rect 45666 66222 45678 66274
rect 50194 66222 50206 66274
rect 50258 66222 50270 66274
rect 54562 66222 54574 66274
rect 54626 66222 54638 66274
rect 54798 66210 54850 66222
rect 54910 66274 54962 66286
rect 54910 66210 54962 66222
rect 55246 66274 55298 66286
rect 55246 66210 55298 66222
rect 56590 66274 56642 66286
rect 56590 66210 56642 66222
rect 56702 66274 56754 66286
rect 56702 66210 56754 66222
rect 57038 66274 57090 66286
rect 57038 66210 57090 66222
rect 57598 66274 57650 66286
rect 75182 66274 75234 66286
rect 78206 66274 78258 66286
rect 115054 66274 115106 66286
rect 58482 66222 58494 66274
rect 58546 66222 58558 66274
rect 61506 66222 61518 66274
rect 61570 66222 61582 66274
rect 62962 66222 62974 66274
rect 63026 66222 63038 66274
rect 71362 66222 71374 66274
rect 71426 66222 71438 66274
rect 75618 66222 75630 66274
rect 75682 66222 75694 66274
rect 114146 66222 114158 66274
rect 114210 66222 114222 66274
rect 57598 66210 57650 66222
rect 75182 66210 75234 66222
rect 78206 66210 78258 66222
rect 115054 66210 115106 66222
rect 115390 66274 115442 66286
rect 115390 66210 115442 66222
rect 117406 66274 117458 66286
rect 117406 66210 117458 66222
rect 52334 66162 52386 66174
rect 1922 66110 1934 66162
rect 1986 66110 1998 66162
rect 52334 66098 52386 66110
rect 52670 66162 52722 66174
rect 52670 66098 52722 66110
rect 54014 66162 54066 66174
rect 54014 66098 54066 66110
rect 58158 66162 58210 66174
rect 58158 66098 58210 66110
rect 61742 66162 61794 66174
rect 77198 66162 77250 66174
rect 113486 66162 113538 66174
rect 117070 66162 117122 66174
rect 75954 66110 75966 66162
rect 76018 66110 76030 66162
rect 78418 66110 78430 66162
rect 78482 66110 78494 66162
rect 78866 66110 78878 66162
rect 78930 66110 78942 66162
rect 115602 66110 115614 66162
rect 115666 66110 115678 66162
rect 116050 66110 116062 66162
rect 116114 66110 116126 66162
rect 61742 66098 61794 66110
rect 77198 66098 77250 66110
rect 113486 66098 113538 66110
rect 117070 66098 117122 66110
rect 117854 66162 117906 66174
rect 117854 66098 117906 66110
rect 45838 66050 45890 66062
rect 45838 65986 45890 65998
rect 50654 66050 50706 66062
rect 50654 65986 50706 65998
rect 51886 66050 51938 66062
rect 51886 65986 51938 65998
rect 53790 66050 53842 66062
rect 53790 65986 53842 65998
rect 55358 66050 55410 66062
rect 55358 65986 55410 65998
rect 56478 66050 56530 66062
rect 56478 65986 56530 65998
rect 57710 66050 57762 66062
rect 57710 65986 57762 65998
rect 62190 66050 62242 66062
rect 62190 65986 62242 65998
rect 66334 66050 66386 66062
rect 66334 65986 66386 65998
rect 66782 66050 66834 66062
rect 66782 65986 66834 65998
rect 67342 66050 67394 66062
rect 67342 65986 67394 65998
rect 69246 66050 69298 66062
rect 69246 65986 69298 65998
rect 81678 66050 81730 66062
rect 81678 65986 81730 65998
rect 114382 66050 114434 66062
rect 114382 65986 114434 65998
rect 1344 65882 118608 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 81278 65882
rect 81330 65830 81382 65882
rect 81434 65830 81486 65882
rect 81538 65830 111998 65882
rect 112050 65830 112102 65882
rect 112154 65830 112206 65882
rect 112258 65830 118608 65882
rect 1344 65796 118608 65830
rect 1822 65714 1874 65726
rect 1822 65650 1874 65662
rect 54686 65714 54738 65726
rect 54686 65650 54738 65662
rect 55022 65714 55074 65726
rect 77422 65714 77474 65726
rect 55570 65662 55582 65714
rect 55634 65662 55646 65714
rect 63298 65662 63310 65714
rect 63362 65662 63374 65714
rect 55022 65650 55074 65662
rect 77422 65650 77474 65662
rect 113934 65714 113986 65726
rect 113934 65650 113986 65662
rect 58494 65602 58546 65614
rect 46722 65550 46734 65602
rect 46786 65550 46798 65602
rect 58494 65538 58546 65550
rect 62302 65602 62354 65614
rect 115266 65550 115278 65602
rect 115330 65550 115342 65602
rect 62302 65538 62354 65550
rect 47966 65490 48018 65502
rect 47506 65438 47518 65490
rect 47570 65438 47582 65490
rect 47966 65426 48018 65438
rect 49534 65490 49586 65502
rect 49534 65426 49586 65438
rect 49982 65490 50034 65502
rect 49982 65426 50034 65438
rect 53342 65490 53394 65502
rect 53342 65426 53394 65438
rect 61518 65490 61570 65502
rect 61518 65426 61570 65438
rect 62414 65490 62466 65502
rect 62414 65426 62466 65438
rect 62526 65490 62578 65502
rect 64654 65490 64706 65502
rect 74622 65490 74674 65502
rect 117854 65490 117906 65502
rect 62962 65438 62974 65490
rect 63026 65438 63038 65490
rect 65650 65438 65662 65490
rect 65714 65438 65726 65490
rect 69122 65438 69134 65490
rect 69186 65438 69198 65490
rect 114482 65438 114494 65490
rect 114546 65438 114558 65490
rect 62526 65426 62578 65438
rect 64654 65426 64706 65438
rect 74622 65426 74674 65438
rect 117854 65426 117906 65438
rect 48750 65378 48802 65390
rect 44594 65326 44606 65378
rect 44658 65326 44670 65378
rect 48750 65314 48802 65326
rect 53790 65378 53842 65390
rect 53790 65314 53842 65326
rect 54238 65378 54290 65390
rect 54238 65314 54290 65326
rect 55918 65378 55970 65390
rect 55918 65314 55970 65326
rect 56142 65378 56194 65390
rect 56142 65314 56194 65326
rect 56590 65378 56642 65390
rect 56590 65314 56642 65326
rect 57486 65378 57538 65390
rect 57486 65314 57538 65326
rect 58046 65378 58098 65390
rect 58046 65314 58098 65326
rect 59838 65378 59890 65390
rect 59838 65314 59890 65326
rect 60958 65378 61010 65390
rect 60958 65314 61010 65326
rect 63198 65378 63250 65390
rect 63198 65314 63250 65326
rect 63534 65378 63586 65390
rect 63534 65314 63586 65326
rect 63870 65378 63922 65390
rect 74174 65378 74226 65390
rect 66434 65326 66446 65378
rect 66498 65326 66510 65378
rect 68562 65326 68574 65378
rect 68626 65326 68638 65378
rect 69906 65326 69918 65378
rect 69970 65326 69982 65378
rect 72034 65326 72046 65378
rect 72098 65326 72110 65378
rect 63870 65314 63922 65326
rect 74174 65314 74226 65326
rect 75070 65378 75122 65390
rect 117394 65326 117406 65378
rect 117458 65326 117470 65378
rect 75070 65314 75122 65326
rect 1344 65098 118608 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 96638 65098
rect 96690 65046 96742 65098
rect 96794 65046 96846 65098
rect 96898 65046 118608 65098
rect 1344 65012 118608 65046
rect 45614 64930 45666 64942
rect 62178 64878 62190 64930
rect 62242 64927 62254 64930
rect 62514 64927 62526 64930
rect 62242 64881 62526 64927
rect 62242 64878 62254 64881
rect 62514 64878 62526 64881
rect 62578 64878 62590 64930
rect 45614 64866 45666 64878
rect 44718 64818 44770 64830
rect 44718 64754 44770 64766
rect 54910 64818 54962 64830
rect 60174 64818 60226 64830
rect 57138 64766 57150 64818
rect 57202 64766 57214 64818
rect 54910 64754 54962 64766
rect 60174 64754 60226 64766
rect 62190 64818 62242 64830
rect 62190 64754 62242 64766
rect 62638 64818 62690 64830
rect 62638 64754 62690 64766
rect 63422 64818 63474 64830
rect 63422 64754 63474 64766
rect 68014 64818 68066 64830
rect 68014 64754 68066 64766
rect 72158 64818 72210 64830
rect 116958 64818 117010 64830
rect 114818 64766 114830 64818
rect 114882 64766 114894 64818
rect 72158 64754 72210 64766
rect 116958 64754 117010 64766
rect 45950 64706 46002 64718
rect 55358 64706 55410 64718
rect 60622 64706 60674 64718
rect 65326 64706 65378 64718
rect 46722 64654 46734 64706
rect 46786 64654 46798 64706
rect 57810 64654 57822 64706
rect 57874 64654 57886 64706
rect 58818 64654 58830 64706
rect 58882 64654 58894 64706
rect 63634 64654 63646 64706
rect 63698 64654 63710 64706
rect 64082 64654 64094 64706
rect 64146 64654 64158 64706
rect 45950 64642 46002 64654
rect 55358 64642 55410 64654
rect 60622 64642 60674 64654
rect 65326 64642 65378 64654
rect 65998 64706 66050 64718
rect 65998 64642 66050 64654
rect 68462 64706 68514 64718
rect 68462 64642 68514 64654
rect 69358 64706 69410 64718
rect 69358 64642 69410 64654
rect 47854 64594 47906 64606
rect 46498 64542 46510 64594
rect 46562 64542 46574 64594
rect 47854 64530 47906 64542
rect 48190 64594 48242 64606
rect 48190 64530 48242 64542
rect 48414 64594 48466 64606
rect 66446 64594 66498 64606
rect 57922 64542 57934 64594
rect 57986 64542 57998 64594
rect 58930 64542 58942 64594
rect 58994 64542 59006 64594
rect 48414 64530 48466 64542
rect 66446 64530 66498 64542
rect 66670 64594 66722 64606
rect 69694 64594 69746 64606
rect 67666 64542 67678 64594
rect 67730 64542 67742 64594
rect 66670 64530 66722 64542
rect 69694 64530 69746 64542
rect 69918 64594 69970 64606
rect 69918 64530 69970 64542
rect 70478 64594 70530 64606
rect 70478 64530 70530 64542
rect 70590 64594 70642 64606
rect 70590 64530 70642 64542
rect 70702 64594 70754 64606
rect 116162 64542 116174 64594
rect 116226 64542 116238 64594
rect 70702 64530 70754 64542
rect 1822 64482 1874 64494
rect 1822 64418 1874 64430
rect 47294 64482 47346 64494
rect 47294 64418 47346 64430
rect 47966 64482 48018 64494
rect 47966 64418 48018 64430
rect 49198 64482 49250 64494
rect 49198 64418 49250 64430
rect 49646 64482 49698 64494
rect 49646 64418 49698 64430
rect 50206 64482 50258 64494
rect 50206 64418 50258 64430
rect 50654 64482 50706 64494
rect 50654 64418 50706 64430
rect 54238 64482 54290 64494
rect 54238 64418 54290 64430
rect 55694 64482 55746 64494
rect 55694 64418 55746 64430
rect 65438 64482 65490 64494
rect 65438 64418 65490 64430
rect 66334 64482 66386 64494
rect 66334 64418 66386 64430
rect 67118 64482 67170 64494
rect 67118 64418 67170 64430
rect 69582 64482 69634 64494
rect 69582 64418 69634 64430
rect 71262 64482 71314 64494
rect 71262 64418 71314 64430
rect 71710 64482 71762 64494
rect 71710 64418 71762 64430
rect 1344 64314 118608 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 81278 64314
rect 81330 64262 81382 64314
rect 81434 64262 81486 64314
rect 81538 64262 111998 64314
rect 112050 64262 112102 64314
rect 112154 64262 112206 64314
rect 112258 64262 118608 64314
rect 1344 64228 118608 64262
rect 53454 64146 53506 64158
rect 53454 64082 53506 64094
rect 54126 64146 54178 64158
rect 54126 64082 54178 64094
rect 56702 64146 56754 64158
rect 56702 64082 56754 64094
rect 58382 64146 58434 64158
rect 58382 64082 58434 64094
rect 63086 64146 63138 64158
rect 63086 64082 63138 64094
rect 65550 64146 65602 64158
rect 65550 64082 65602 64094
rect 66558 64146 66610 64158
rect 66558 64082 66610 64094
rect 68126 64146 68178 64158
rect 68126 64082 68178 64094
rect 68686 64146 68738 64158
rect 68686 64082 68738 64094
rect 70702 64146 70754 64158
rect 70702 64082 70754 64094
rect 49646 64034 49698 64046
rect 1922 63982 1934 64034
rect 1986 63982 1998 64034
rect 47954 63982 47966 64034
rect 48018 63982 48030 64034
rect 49646 63970 49698 63982
rect 62750 64034 62802 64046
rect 62750 63970 62802 63982
rect 65662 64034 65714 64046
rect 65662 63970 65714 63982
rect 67342 64034 67394 64046
rect 67342 63970 67394 63982
rect 51214 63922 51266 63934
rect 55806 63922 55858 63934
rect 48626 63870 48638 63922
rect 48690 63870 48702 63922
rect 50754 63870 50766 63922
rect 50818 63870 50830 63922
rect 55346 63870 55358 63922
rect 55410 63870 55422 63922
rect 51214 63858 51266 63870
rect 55806 63858 55858 63870
rect 57598 63922 57650 63934
rect 64766 63922 64818 63934
rect 59042 63870 59054 63922
rect 59106 63870 59118 63922
rect 59826 63870 59838 63922
rect 59890 63870 59902 63922
rect 64194 63870 64206 63922
rect 64258 63870 64270 63922
rect 57598 63858 57650 63870
rect 64766 63858 64818 63870
rect 65326 63922 65378 63934
rect 69470 63922 69522 63934
rect 71150 63922 71202 63934
rect 67666 63870 67678 63922
rect 67730 63870 67742 63922
rect 70466 63870 70478 63922
rect 70530 63870 70542 63922
rect 65326 63858 65378 63870
rect 69470 63858 69522 63870
rect 71150 63858 71202 63870
rect 50430 63810 50482 63822
rect 3266 63758 3278 63810
rect 3330 63758 3342 63810
rect 45826 63758 45838 63810
rect 45890 63758 45902 63810
rect 49522 63758 49534 63810
rect 49586 63758 49598 63810
rect 50430 63746 50482 63758
rect 50542 63810 50594 63822
rect 50542 63746 50594 63758
rect 54238 63810 54290 63822
rect 54238 63746 54290 63758
rect 54910 63810 54962 63822
rect 63646 63810 63698 63822
rect 58482 63758 58494 63810
rect 58546 63758 58558 63810
rect 61954 63758 61966 63810
rect 62018 63758 62030 63810
rect 54910 63746 54962 63758
rect 63646 63746 63698 63758
rect 63758 63810 63810 63822
rect 63758 63746 63810 63758
rect 66222 63810 66274 63822
rect 66222 63746 66274 63758
rect 67454 63810 67506 63822
rect 67454 63746 67506 63758
rect 69022 63810 69074 63822
rect 69022 63746 69074 63758
rect 49870 63698 49922 63710
rect 49870 63634 49922 63646
rect 54350 63698 54402 63710
rect 54350 63634 54402 63646
rect 58158 63698 58210 63710
rect 58158 63634 58210 63646
rect 63982 63698 64034 63710
rect 63982 63634 64034 63646
rect 1344 63530 118608 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 96638 63530
rect 96690 63478 96742 63530
rect 96794 63478 96846 63530
rect 96898 63478 118608 63530
rect 1344 63444 118608 63478
rect 63198 63362 63250 63374
rect 51762 63310 51774 63362
rect 51826 63359 51838 63362
rect 51986 63359 51998 63362
rect 51826 63313 51998 63359
rect 51826 63310 51838 63313
rect 51986 63310 51998 63313
rect 52050 63310 52062 63362
rect 63198 63298 63250 63310
rect 51998 63250 52050 63262
rect 56366 63250 56418 63262
rect 3266 63198 3278 63250
rect 3330 63198 3342 63250
rect 48626 63198 48638 63250
rect 48690 63198 48702 63250
rect 54226 63198 54238 63250
rect 54290 63198 54302 63250
rect 51998 63186 52050 63198
rect 56366 63186 56418 63198
rect 57374 63250 57426 63262
rect 57374 63186 57426 63198
rect 57822 63250 57874 63262
rect 57822 63186 57874 63198
rect 58270 63250 58322 63262
rect 68014 63250 68066 63262
rect 62850 63198 62862 63250
rect 62914 63198 62926 63250
rect 58270 63186 58322 63198
rect 68014 63186 68066 63198
rect 70142 63250 70194 63262
rect 74498 63198 74510 63250
rect 74562 63198 74574 63250
rect 114818 63198 114830 63250
rect 114882 63198 114894 63250
rect 70142 63186 70194 63198
rect 58606 63138 58658 63150
rect 47618 63086 47630 63138
rect 47682 63086 47694 63138
rect 51538 63086 51550 63138
rect 51602 63086 51614 63138
rect 53554 63086 53566 63138
rect 53618 63086 53630 63138
rect 58606 63074 58658 63086
rect 58942 63138 58994 63150
rect 59614 63138 59666 63150
rect 59154 63086 59166 63138
rect 59218 63086 59230 63138
rect 58942 63074 58994 63086
rect 59614 63074 59666 63086
rect 65438 63138 65490 63150
rect 65762 63086 65774 63138
rect 65826 63086 65838 63138
rect 71586 63086 71598 63138
rect 71650 63086 71662 63138
rect 65438 63074 65490 63086
rect 48078 63026 48130 63038
rect 58494 63026 58546 63038
rect 1922 62974 1934 63026
rect 1986 62974 1998 63026
rect 50754 62974 50766 63026
rect 50818 62974 50830 63026
rect 48078 62962 48130 62974
rect 58494 62962 58546 62974
rect 61406 63026 61458 63038
rect 61406 62962 61458 62974
rect 62078 63026 62130 63038
rect 62078 62962 62130 62974
rect 62190 63026 62242 63038
rect 64318 63026 64370 63038
rect 62402 62974 62414 63026
rect 62466 63023 62478 63026
rect 62738 63023 62750 63026
rect 62466 62977 62750 63023
rect 62466 62974 62478 62977
rect 62738 62974 62750 62977
rect 62802 62974 62814 63026
rect 62190 62962 62242 62974
rect 64318 62962 64370 62974
rect 66334 63026 66386 63038
rect 66334 62962 66386 62974
rect 69358 63026 69410 63038
rect 72370 62974 72382 63026
rect 72434 62974 72446 63026
rect 116162 62974 116174 63026
rect 116226 62974 116238 63026
rect 69358 62962 69410 62974
rect 58158 62914 58210 62926
rect 58158 62850 58210 62862
rect 61854 62914 61906 62926
rect 61854 62850 61906 62862
rect 62974 62914 63026 62926
rect 68462 62914 68514 62926
rect 63858 62862 63870 62914
rect 63922 62862 63934 62914
rect 62974 62850 63026 62862
rect 68462 62850 68514 62862
rect 69470 62914 69522 62926
rect 69470 62850 69522 62862
rect 71038 62914 71090 62926
rect 71038 62850 71090 62862
rect 74958 62914 75010 62926
rect 74958 62850 75010 62862
rect 117070 62914 117122 62926
rect 117070 62850 117122 62862
rect 1344 62746 118608 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 81278 62746
rect 81330 62694 81382 62746
rect 81434 62694 81486 62746
rect 81538 62694 111998 62746
rect 112050 62694 112102 62746
rect 112154 62694 112206 62746
rect 112258 62694 118608 62746
rect 1344 62660 118608 62694
rect 1822 62578 1874 62590
rect 1822 62514 1874 62526
rect 50318 62578 50370 62590
rect 50318 62514 50370 62526
rect 54686 62578 54738 62590
rect 54686 62514 54738 62526
rect 55246 62578 55298 62590
rect 55246 62514 55298 62526
rect 56254 62578 56306 62590
rect 56254 62514 56306 62526
rect 63086 62578 63138 62590
rect 63086 62514 63138 62526
rect 63758 62578 63810 62590
rect 63758 62514 63810 62526
rect 64654 62578 64706 62590
rect 64654 62514 64706 62526
rect 70030 62578 70082 62590
rect 70030 62514 70082 62526
rect 72046 62578 72098 62590
rect 72046 62514 72098 62526
rect 45838 62466 45890 62478
rect 45838 62402 45890 62414
rect 49534 62466 49586 62478
rect 49534 62402 49586 62414
rect 50094 62466 50146 62478
rect 50094 62402 50146 62414
rect 55134 62466 55186 62478
rect 55134 62402 55186 62414
rect 56702 62466 56754 62478
rect 56702 62402 56754 62414
rect 58494 62466 58546 62478
rect 58494 62402 58546 62414
rect 58942 62466 58994 62478
rect 58942 62402 58994 62414
rect 73390 62466 73442 62478
rect 73390 62402 73442 62414
rect 74174 62466 74226 62478
rect 74174 62402 74226 62414
rect 45502 62354 45554 62366
rect 45502 62290 45554 62302
rect 50430 62354 50482 62366
rect 50430 62290 50482 62302
rect 50542 62354 50594 62366
rect 50542 62290 50594 62302
rect 51102 62354 51154 62366
rect 51102 62290 51154 62302
rect 52894 62354 52946 62366
rect 55022 62354 55074 62366
rect 63646 62354 63698 62366
rect 54450 62302 54462 62354
rect 54514 62302 54526 62354
rect 58034 62302 58046 62354
rect 58098 62302 58110 62354
rect 61842 62302 61854 62354
rect 61906 62302 61918 62354
rect 62514 62302 62526 62354
rect 62578 62302 62590 62354
rect 52894 62290 52946 62302
rect 55022 62290 55074 62302
rect 63646 62290 63698 62302
rect 63870 62354 63922 62366
rect 63870 62290 63922 62302
rect 64094 62354 64146 62366
rect 65662 62354 65714 62366
rect 71710 62354 71762 62366
rect 65426 62302 65438 62354
rect 65490 62302 65502 62354
rect 66770 62302 66782 62354
rect 66834 62302 66846 62354
rect 64094 62290 64146 62302
rect 65662 62290 65714 62302
rect 71710 62290 71762 62302
rect 72046 62354 72098 62366
rect 72046 62290 72098 62302
rect 72382 62354 72434 62366
rect 72382 62290 72434 62302
rect 73502 62354 73554 62366
rect 74734 62354 74786 62366
rect 73714 62302 73726 62354
rect 73778 62302 73790 62354
rect 73502 62290 73554 62302
rect 74734 62290 74786 62302
rect 48302 62242 48354 62254
rect 48302 62178 48354 62190
rect 53342 62242 53394 62254
rect 53342 62178 53394 62190
rect 53790 62242 53842 62254
rect 53790 62178 53842 62190
rect 55470 62242 55522 62254
rect 55470 62178 55522 62190
rect 55806 62242 55858 62254
rect 70478 62242 70530 62254
rect 57586 62190 57598 62242
rect 57650 62190 57662 62242
rect 59714 62190 59726 62242
rect 59778 62190 59790 62242
rect 67442 62190 67454 62242
rect 67506 62190 67518 62242
rect 69570 62190 69582 62242
rect 69634 62190 69646 62242
rect 55806 62178 55858 62190
rect 70478 62178 70530 62190
rect 70926 62242 70978 62254
rect 70926 62178 70978 62190
rect 53902 62130 53954 62142
rect 53902 62066 53954 62078
rect 65774 62130 65826 62142
rect 65774 62066 65826 62078
rect 1344 61962 118608 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 96638 61962
rect 96690 61910 96742 61962
rect 96794 61910 96846 61962
rect 96898 61910 118608 61962
rect 1344 61876 118608 61910
rect 54014 61794 54066 61806
rect 55906 61742 55918 61794
rect 55970 61791 55982 61794
rect 56466 61791 56478 61794
rect 55970 61745 56478 61791
rect 55970 61742 55982 61745
rect 56466 61742 56478 61745
rect 56530 61742 56542 61794
rect 57810 61742 57822 61794
rect 57874 61791 57886 61794
rect 58818 61791 58830 61794
rect 57874 61745 58830 61791
rect 57874 61742 57886 61745
rect 58818 61742 58830 61745
rect 58882 61742 58894 61794
rect 54014 61730 54066 61742
rect 3614 61682 3666 61694
rect 48862 61682 48914 61694
rect 46274 61630 46286 61682
rect 46338 61630 46350 61682
rect 48402 61630 48414 61682
rect 48466 61630 48478 61682
rect 3614 61618 3666 61630
rect 48862 61618 48914 61630
rect 49310 61682 49362 61694
rect 49310 61618 49362 61630
rect 51214 61682 51266 61694
rect 51214 61618 51266 61630
rect 53566 61682 53618 61694
rect 53566 61618 53618 61630
rect 55582 61682 55634 61694
rect 55582 61618 55634 61630
rect 55918 61682 55970 61694
rect 55918 61618 55970 61630
rect 59278 61682 59330 61694
rect 59278 61618 59330 61630
rect 59726 61682 59778 61694
rect 68350 61682 68402 61694
rect 62514 61630 62526 61682
rect 62578 61630 62590 61682
rect 59726 61618 59778 61630
rect 68350 61618 68402 61630
rect 70814 61682 70866 61694
rect 74498 61630 74510 61682
rect 74562 61630 74574 61682
rect 80434 61630 80446 61682
rect 80498 61630 80510 61682
rect 114818 61630 114830 61682
rect 114882 61630 114894 61682
rect 70814 61618 70866 61630
rect 67454 61570 67506 61582
rect 69470 61570 69522 61582
rect 3042 61518 3054 61570
rect 3106 61518 3118 61570
rect 45602 61518 45614 61570
rect 45666 61518 45678 61570
rect 66658 61518 66670 61570
rect 66722 61518 66734 61570
rect 67890 61518 67902 61570
rect 67954 61518 67966 61570
rect 67454 61506 67506 61518
rect 69470 61506 69522 61518
rect 69918 61570 69970 61582
rect 83022 61570 83074 61582
rect 71698 61518 71710 61570
rect 71762 61518 71774 61570
rect 81106 61518 81118 61570
rect 81170 61518 81182 61570
rect 69918 61506 69970 61518
rect 83022 61506 83074 61518
rect 54350 61458 54402 61470
rect 1922 61406 1934 61458
rect 1986 61406 1998 61458
rect 54350 61394 54402 61406
rect 67566 61458 67618 61470
rect 67566 61394 67618 61406
rect 70926 61458 70978 61470
rect 72370 61406 72382 61458
rect 72434 61406 72446 61458
rect 116162 61406 116174 61458
rect 116226 61406 116238 61458
rect 70926 61394 70978 61406
rect 50878 61346 50930 61358
rect 50878 61282 50930 61294
rect 52222 61346 52274 61358
rect 52222 61282 52274 61294
rect 52670 61346 52722 61358
rect 52670 61282 52722 61294
rect 54126 61346 54178 61358
rect 54126 61282 54178 61294
rect 55022 61346 55074 61358
rect 55022 61282 55074 61294
rect 56366 61346 56418 61358
rect 56366 61282 56418 61294
rect 56814 61346 56866 61358
rect 56814 61282 56866 61294
rect 57598 61346 57650 61358
rect 57598 61282 57650 61294
rect 58046 61346 58098 61358
rect 58046 61282 58098 61294
rect 58494 61346 58546 61358
rect 58494 61282 58546 61294
rect 58942 61346 58994 61358
rect 58942 61282 58994 61294
rect 67342 61346 67394 61358
rect 67342 61282 67394 61294
rect 67678 61346 67730 61358
rect 67678 61282 67730 61294
rect 70030 61346 70082 61358
rect 70030 61282 70082 61294
rect 70142 61346 70194 61358
rect 70142 61282 70194 61294
rect 74958 61346 75010 61358
rect 74958 61282 75010 61294
rect 117070 61346 117122 61358
rect 117070 61282 117122 61294
rect 1344 61178 118608 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 81278 61178
rect 81330 61126 81382 61178
rect 81434 61126 81486 61178
rect 81538 61126 111998 61178
rect 112050 61126 112102 61178
rect 112154 61126 112206 61178
rect 112258 61126 118608 61178
rect 1344 61092 118608 61126
rect 45726 61010 45778 61022
rect 45726 60946 45778 60958
rect 52670 61010 52722 61022
rect 52670 60946 52722 60958
rect 59390 61010 59442 61022
rect 59390 60946 59442 60958
rect 60286 61010 60338 61022
rect 60286 60946 60338 60958
rect 61518 61010 61570 61022
rect 61518 60946 61570 60958
rect 67678 61010 67730 61022
rect 67678 60946 67730 60958
rect 68574 61010 68626 61022
rect 68574 60946 68626 60958
rect 69470 61010 69522 61022
rect 69470 60946 69522 60958
rect 71934 61010 71986 61022
rect 71934 60946 71986 60958
rect 73614 61010 73666 61022
rect 73614 60946 73666 60958
rect 74286 61010 74338 61022
rect 74286 60946 74338 60958
rect 56366 60898 56418 60910
rect 46610 60846 46622 60898
rect 46674 60846 46686 60898
rect 56366 60834 56418 60846
rect 58382 60898 58434 60910
rect 58382 60834 58434 60846
rect 59614 60898 59666 60910
rect 59614 60834 59666 60846
rect 59838 60898 59890 60910
rect 59838 60834 59890 60846
rect 61742 60898 61794 60910
rect 61742 60834 61794 60846
rect 65662 60898 65714 60910
rect 65662 60834 65714 60846
rect 67454 60898 67506 60910
rect 67454 60834 67506 60846
rect 68014 60898 68066 60910
rect 68014 60834 68066 60846
rect 70366 60898 70418 60910
rect 70366 60834 70418 60846
rect 70926 60898 70978 60910
rect 116274 60846 116286 60898
rect 116338 60846 116350 60898
rect 70926 60834 70978 60846
rect 46062 60786 46114 60798
rect 53566 60786 53618 60798
rect 55134 60786 55186 60798
rect 58494 60786 58546 60798
rect 59502 60786 59554 60798
rect 46498 60734 46510 60786
rect 46562 60734 46574 60786
rect 47730 60734 47742 60786
rect 47794 60734 47806 60786
rect 50194 60734 50206 60786
rect 50258 60734 50270 60786
rect 54002 60734 54014 60786
rect 54066 60734 54078 60786
rect 56018 60734 56030 60786
rect 56082 60734 56094 60786
rect 59154 60734 59166 60786
rect 59218 60734 59230 60786
rect 46062 60722 46114 60734
rect 53566 60722 53618 60734
rect 55134 60722 55186 60734
rect 58494 60722 58546 60734
rect 59502 60722 59554 60734
rect 61294 60786 61346 60798
rect 61294 60722 61346 60734
rect 61966 60786 62018 60798
rect 61966 60722 62018 60734
rect 62414 60786 62466 60798
rect 67790 60786 67842 60798
rect 63522 60734 63534 60786
rect 63586 60734 63598 60786
rect 62414 60722 62466 60734
rect 67790 60722 67842 60734
rect 69582 60786 69634 60798
rect 69582 60722 69634 60734
rect 69806 60786 69858 60798
rect 69806 60722 69858 60734
rect 70254 60786 70306 60798
rect 70254 60722 70306 60734
rect 71598 60786 71650 60798
rect 71598 60722 71650 60734
rect 71934 60786 71986 60798
rect 71934 60722 71986 60734
rect 72270 60786 72322 60798
rect 72270 60722 72322 60734
rect 1822 60674 1874 60686
rect 49534 60674 49586 60686
rect 50990 60674 51042 60686
rect 48178 60622 48190 60674
rect 48242 60622 48254 60674
rect 50306 60622 50318 60674
rect 50370 60622 50382 60674
rect 1822 60610 1874 60622
rect 49534 60610 49586 60622
rect 50990 60610 51042 60622
rect 51550 60674 51602 60686
rect 51550 60610 51602 60622
rect 52222 60674 52274 60686
rect 52222 60610 52274 60622
rect 53006 60674 53058 60686
rect 53006 60610 53058 60622
rect 57710 60674 57762 60686
rect 57710 60610 57762 60622
rect 60734 60674 60786 60686
rect 60734 60610 60786 60622
rect 62974 60674 63026 60686
rect 64430 60674 64482 60686
rect 63746 60622 63758 60674
rect 63810 60622 63822 60674
rect 62974 60610 63026 60622
rect 64430 60610 64482 60622
rect 66222 60674 66274 60686
rect 66222 60610 66274 60622
rect 66670 60674 66722 60686
rect 66670 60610 66722 60622
rect 68686 60674 68738 60686
rect 68686 60610 68738 60622
rect 71038 60674 71090 60686
rect 116846 60674 116898 60686
rect 73602 60622 73614 60674
rect 73666 60622 73678 60674
rect 114930 60622 114942 60674
rect 114994 60622 115006 60674
rect 71038 60610 71090 60622
rect 116846 60610 116898 60622
rect 54014 60562 54066 60574
rect 54014 60498 54066 60510
rect 54350 60562 54402 60574
rect 54350 60498 54402 60510
rect 55022 60562 55074 60574
rect 55022 60498 55074 60510
rect 55358 60562 55410 60574
rect 55358 60498 55410 60510
rect 55470 60562 55522 60574
rect 55470 60498 55522 60510
rect 56030 60562 56082 60574
rect 56030 60498 56082 60510
rect 58606 60562 58658 60574
rect 58606 60498 58658 60510
rect 65438 60562 65490 60574
rect 65438 60498 65490 60510
rect 65774 60562 65826 60574
rect 73390 60562 73442 60574
rect 66210 60510 66222 60562
rect 66274 60559 66286 60562
rect 66770 60559 66782 60562
rect 66274 60513 66782 60559
rect 66274 60510 66286 60513
rect 66770 60510 66782 60513
rect 66834 60510 66846 60562
rect 65774 60498 65826 60510
rect 73390 60498 73442 60510
rect 1344 60394 118608 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 96638 60394
rect 96690 60342 96742 60394
rect 96794 60342 96846 60394
rect 96898 60342 118608 60394
rect 1344 60308 118608 60342
rect 55358 60226 55410 60238
rect 51202 60174 51214 60226
rect 51266 60223 51278 60226
rect 51874 60223 51886 60226
rect 51266 60177 51886 60223
rect 51266 60174 51278 60177
rect 51874 60174 51886 60177
rect 51938 60174 51950 60226
rect 55358 60162 55410 60174
rect 58718 60226 58770 60238
rect 58718 60162 58770 60174
rect 59502 60226 59554 60238
rect 59502 60162 59554 60174
rect 59950 60226 60002 60238
rect 68014 60226 68066 60238
rect 62290 60174 62302 60226
rect 62354 60223 62366 60226
rect 63074 60223 63086 60226
rect 62354 60177 63086 60223
rect 62354 60174 62366 60177
rect 63074 60174 63086 60177
rect 63138 60174 63150 60226
rect 59950 60162 60002 60174
rect 68014 60162 68066 60174
rect 69918 60226 69970 60238
rect 69918 60162 69970 60174
rect 47070 60114 47122 60126
rect 3266 60062 3278 60114
rect 3330 60062 3342 60114
rect 47070 60050 47122 60062
rect 47966 60114 48018 60126
rect 47966 60050 48018 60062
rect 49198 60114 49250 60126
rect 49198 60050 49250 60062
rect 49646 60114 49698 60126
rect 61294 60114 61346 60126
rect 53890 60062 53902 60114
rect 53954 60062 53966 60114
rect 56466 60062 56478 60114
rect 56530 60062 56542 60114
rect 58482 60062 58494 60114
rect 58546 60062 58558 60114
rect 49646 60050 49698 60062
rect 61294 60050 61346 60062
rect 61854 60114 61906 60126
rect 61854 60050 61906 60062
rect 62302 60114 62354 60126
rect 67006 60114 67058 60126
rect 63522 60062 63534 60114
rect 63586 60062 63598 60114
rect 65762 60062 65774 60114
rect 65826 60062 65838 60114
rect 62302 60050 62354 60062
rect 67006 60050 67058 60062
rect 67454 60114 67506 60126
rect 67454 60050 67506 60062
rect 70478 60114 70530 60126
rect 70478 60050 70530 60062
rect 71822 60114 71874 60126
rect 71822 60050 71874 60062
rect 48750 60002 48802 60014
rect 50206 60002 50258 60014
rect 49746 59950 49758 60002
rect 49810 59950 49822 60002
rect 48750 59938 48802 59950
rect 50206 59938 50258 59950
rect 50318 60002 50370 60014
rect 50318 59938 50370 59950
rect 50430 60002 50482 60014
rect 50430 59938 50482 59950
rect 51886 60002 51938 60014
rect 55134 60002 55186 60014
rect 55918 60002 55970 60014
rect 57822 60002 57874 60014
rect 53554 59950 53566 60002
rect 53618 59950 53630 60002
rect 55570 59950 55582 60002
rect 55634 59950 55646 60002
rect 57026 59950 57038 60002
rect 57090 59950 57102 60002
rect 51886 59938 51938 59950
rect 55134 59938 55186 59950
rect 55918 59938 55970 59950
rect 57822 59938 57874 59950
rect 59390 60002 59442 60014
rect 59390 59938 59442 59950
rect 59726 60002 59778 60014
rect 68686 60002 68738 60014
rect 66546 59950 66558 60002
rect 66610 59950 66622 60002
rect 59726 59938 59778 59950
rect 68686 59938 68738 59950
rect 69358 60002 69410 60014
rect 69358 59938 69410 59950
rect 71374 60002 71426 60014
rect 71374 59938 71426 59950
rect 47406 59890 47458 59902
rect 1922 59838 1934 59890
rect 1986 59838 1998 59890
rect 47406 59826 47458 59838
rect 52782 59890 52834 59902
rect 52782 59826 52834 59838
rect 54910 59890 54962 59902
rect 57710 59890 57762 59902
rect 70030 59890 70082 59902
rect 56690 59838 56702 59890
rect 56754 59838 56766 59890
rect 62962 59838 62974 59890
rect 63026 59887 63038 59890
rect 63298 59887 63310 59890
rect 63026 59841 63310 59887
rect 63026 59838 63038 59841
rect 63298 59838 63310 59841
rect 63362 59838 63374 59890
rect 54910 59826 54962 59838
rect 57710 59826 57762 59838
rect 70030 59826 70082 59838
rect 46510 59778 46562 59790
rect 46510 59714 46562 59726
rect 48302 59778 48354 59790
rect 48302 59714 48354 59726
rect 49534 59778 49586 59790
rect 49534 59714 49586 59726
rect 51326 59778 51378 59790
rect 51326 59714 51378 59726
rect 52334 59778 52386 59790
rect 52334 59714 52386 59726
rect 54798 59778 54850 59790
rect 54798 59714 54850 59726
rect 57486 59778 57538 59790
rect 57486 59714 57538 59726
rect 58494 59778 58546 59790
rect 58494 59714 58546 59726
rect 59390 59778 59442 59790
rect 59390 59714 59442 59726
rect 60510 59778 60562 59790
rect 60510 59714 60562 59726
rect 62862 59778 62914 59790
rect 62862 59714 62914 59726
rect 68126 59778 68178 59790
rect 68126 59714 68178 59726
rect 68350 59778 68402 59790
rect 68350 59714 68402 59726
rect 69582 59778 69634 59790
rect 69582 59714 69634 59726
rect 69806 59778 69858 59790
rect 69806 59714 69858 59726
rect 70926 59778 70978 59790
rect 70926 59714 70978 59726
rect 73054 59778 73106 59790
rect 115278 59778 115330 59790
rect 114930 59726 114942 59778
rect 114994 59726 115006 59778
rect 73054 59714 73106 59726
rect 115278 59714 115330 59726
rect 115838 59778 115890 59790
rect 115838 59714 115890 59726
rect 1344 59610 118608 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 81278 59610
rect 81330 59558 81382 59610
rect 81434 59558 81486 59610
rect 81538 59558 111998 59610
rect 112050 59558 112102 59610
rect 112154 59558 112206 59610
rect 112258 59558 118608 59610
rect 1344 59524 118608 59558
rect 57822 59442 57874 59454
rect 55010 59390 55022 59442
rect 55074 59390 55086 59442
rect 57822 59378 57874 59390
rect 59950 59442 60002 59454
rect 59950 59378 60002 59390
rect 60958 59442 61010 59454
rect 60958 59378 61010 59390
rect 62862 59442 62914 59454
rect 62862 59378 62914 59390
rect 63646 59442 63698 59454
rect 63646 59378 63698 59390
rect 64318 59442 64370 59454
rect 64318 59378 64370 59390
rect 66782 59442 66834 59454
rect 66782 59378 66834 59390
rect 67566 59442 67618 59454
rect 67566 59378 67618 59390
rect 68910 59442 68962 59454
rect 68910 59378 68962 59390
rect 69358 59442 69410 59454
rect 69358 59378 69410 59390
rect 69694 59442 69746 59454
rect 69694 59378 69746 59390
rect 69918 59442 69970 59454
rect 69918 59378 69970 59390
rect 72046 59442 72098 59454
rect 72046 59378 72098 59390
rect 49534 59330 49586 59342
rect 1922 59278 1934 59330
rect 1986 59278 1998 59330
rect 49534 59266 49586 59278
rect 49758 59330 49810 59342
rect 55582 59330 55634 59342
rect 52882 59278 52894 59330
rect 52946 59278 52958 59330
rect 49758 59266 49810 59278
rect 55582 59266 55634 59278
rect 57598 59330 57650 59342
rect 57598 59266 57650 59278
rect 58494 59330 58546 59342
rect 58494 59266 58546 59278
rect 59054 59330 59106 59342
rect 59054 59266 59106 59278
rect 63310 59330 63362 59342
rect 63310 59266 63362 59278
rect 66110 59330 66162 59342
rect 66110 59266 66162 59278
rect 48750 59218 48802 59230
rect 55918 59218 55970 59230
rect 53554 59166 53566 59218
rect 53618 59166 53630 59218
rect 48750 59154 48802 59166
rect 55918 59154 55970 59166
rect 56366 59218 56418 59230
rect 56366 59154 56418 59166
rect 57486 59218 57538 59230
rect 57486 59154 57538 59166
rect 58718 59218 58770 59230
rect 58718 59154 58770 59166
rect 59614 59218 59666 59230
rect 59614 59154 59666 59166
rect 59950 59218 60002 59230
rect 59950 59154 60002 59166
rect 60286 59218 60338 59230
rect 62078 59218 62130 59230
rect 61170 59166 61182 59218
rect 61234 59166 61246 59218
rect 60286 59154 60338 59166
rect 62078 59154 62130 59166
rect 62750 59218 62802 59230
rect 69470 59218 69522 59230
rect 63074 59166 63086 59218
rect 63138 59166 63150 59218
rect 62750 59154 62802 59166
rect 69470 59154 69522 59166
rect 70142 59218 70194 59230
rect 70142 59154 70194 59166
rect 70590 59218 70642 59230
rect 70590 59154 70642 59166
rect 49646 59106 49698 59118
rect 54462 59106 54514 59118
rect 3266 59054 3278 59106
rect 3330 59054 3342 59106
rect 50754 59054 50766 59106
rect 50818 59054 50830 59106
rect 49646 59042 49698 59054
rect 54462 59042 54514 59054
rect 58942 59106 58994 59118
rect 58942 59042 58994 59054
rect 61630 59106 61682 59118
rect 61630 59042 61682 59054
rect 63534 59106 63586 59118
rect 63534 59042 63586 59054
rect 63982 59106 64034 59118
rect 63982 59042 64034 59054
rect 65326 59106 65378 59118
rect 65326 59042 65378 59054
rect 65886 59106 65938 59118
rect 67118 59106 67170 59118
rect 66210 59054 66222 59106
rect 66274 59054 66286 59106
rect 65886 59042 65938 59054
rect 67118 59042 67170 59054
rect 68014 59106 68066 59118
rect 68014 59042 68066 59054
rect 68462 59106 68514 59118
rect 68462 59042 68514 59054
rect 71038 59106 71090 59118
rect 71038 59042 71090 59054
rect 71486 59106 71538 59118
rect 71486 59042 71538 59054
rect 54686 58994 54738 59006
rect 54686 58930 54738 58942
rect 60846 58994 60898 59006
rect 60846 58930 60898 58942
rect 1344 58826 118608 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 96638 58826
rect 96690 58774 96742 58826
rect 96794 58774 96846 58826
rect 96898 58774 118608 58826
rect 1344 58740 118608 58774
rect 54574 58658 54626 58670
rect 54574 58594 54626 58606
rect 56814 58658 56866 58670
rect 56814 58594 56866 58606
rect 59390 58658 59442 58670
rect 59390 58594 59442 58606
rect 59614 58658 59666 58670
rect 59614 58594 59666 58606
rect 62190 58658 62242 58670
rect 62190 58594 62242 58606
rect 62526 58658 62578 58670
rect 62526 58594 62578 58606
rect 63982 58658 64034 58670
rect 64194 58606 64206 58658
rect 64258 58655 64270 58658
rect 65314 58655 65326 58658
rect 64258 58609 65326 58655
rect 64258 58606 64270 58609
rect 65314 58606 65326 58609
rect 65378 58606 65390 58658
rect 67554 58606 67566 58658
rect 67618 58655 67630 58658
rect 68114 58655 68126 58658
rect 67618 58609 68126 58655
rect 67618 58606 67630 58609
rect 68114 58606 68126 58609
rect 68178 58655 68190 58658
rect 68338 58655 68350 58658
rect 68178 58609 68350 58655
rect 68178 58606 68190 58609
rect 68338 58606 68350 58609
rect 68402 58606 68414 58658
rect 63982 58594 64034 58606
rect 1822 58546 1874 58558
rect 52222 58546 52274 58558
rect 49074 58494 49086 58546
rect 49138 58494 49150 58546
rect 1822 58482 1874 58494
rect 52222 58482 52274 58494
rect 52782 58546 52834 58558
rect 63086 58546 63138 58558
rect 67678 58546 67730 58558
rect 56018 58494 56030 58546
rect 56082 58494 56094 58546
rect 63634 58494 63646 58546
rect 63698 58494 63710 58546
rect 52782 58482 52834 58494
rect 63086 58482 63138 58494
rect 67678 58482 67730 58494
rect 68126 58546 68178 58558
rect 68126 58482 68178 58494
rect 68574 58546 68626 58558
rect 68574 58482 68626 58494
rect 69358 58546 69410 58558
rect 69358 58482 69410 58494
rect 70926 58546 70978 58558
rect 114818 58494 114830 58546
rect 114882 58494 114894 58546
rect 70926 58482 70978 58494
rect 55806 58434 55858 58446
rect 58046 58434 58098 58446
rect 48402 58382 48414 58434
rect 48466 58382 48478 58434
rect 56242 58382 56254 58434
rect 56306 58382 56318 58434
rect 55806 58370 55858 58382
rect 58046 58370 58098 58382
rect 58270 58434 58322 58446
rect 59166 58434 59218 58446
rect 58930 58382 58942 58434
rect 58994 58382 59006 58434
rect 58270 58370 58322 58382
rect 59166 58370 59218 58382
rect 67230 58434 67282 58446
rect 67230 58370 67282 58382
rect 69582 58434 69634 58446
rect 70702 58434 70754 58446
rect 70018 58382 70030 58434
rect 70082 58382 70094 58434
rect 69582 58370 69634 58382
rect 70702 58370 70754 58382
rect 53454 58322 53506 58334
rect 53454 58258 53506 58270
rect 53790 58322 53842 58334
rect 53790 58258 53842 58270
rect 54462 58322 54514 58334
rect 54462 58258 54514 58270
rect 55582 58322 55634 58334
rect 55582 58258 55634 58270
rect 56030 58322 56082 58334
rect 56030 58258 56082 58270
rect 57822 58322 57874 58334
rect 57822 58258 57874 58270
rect 58382 58322 58434 58334
rect 58382 58258 58434 58270
rect 63758 58322 63810 58334
rect 63758 58258 63810 58270
rect 64878 58322 64930 58334
rect 64878 58258 64930 58270
rect 65774 58322 65826 58334
rect 69794 58270 69806 58322
rect 69858 58270 69870 58322
rect 116162 58270 116174 58322
rect 116226 58270 116238 58322
rect 65774 58258 65826 58270
rect 54574 58210 54626 58222
rect 51314 58158 51326 58210
rect 51378 58158 51390 58210
rect 54574 58146 54626 58158
rect 56926 58210 56978 58222
rect 56926 58146 56978 58158
rect 57038 58210 57090 58222
rect 57038 58146 57090 58158
rect 59054 58210 59106 58222
rect 59054 58146 59106 58158
rect 60398 58210 60450 58222
rect 60398 58146 60450 58158
rect 61630 58210 61682 58222
rect 61630 58146 61682 58158
rect 62414 58210 62466 58222
rect 62414 58146 62466 58158
rect 64542 58210 64594 58222
rect 64542 58146 64594 58158
rect 65326 58210 65378 58222
rect 65326 58146 65378 58158
rect 66222 58210 66274 58222
rect 66222 58146 66274 58158
rect 70366 58210 70418 58222
rect 70366 58146 70418 58158
rect 71038 58210 71090 58222
rect 71038 58146 71090 58158
rect 71262 58210 71314 58222
rect 71262 58146 71314 58158
rect 71710 58210 71762 58222
rect 71710 58146 71762 58158
rect 117070 58210 117122 58222
rect 117070 58146 117122 58158
rect 1344 58042 118608 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 81278 58042
rect 81330 57990 81382 58042
rect 81434 57990 81486 58042
rect 81538 57990 111998 58042
rect 112050 57990 112102 58042
rect 112154 57990 112206 58042
rect 112258 57990 118608 58042
rect 1344 57956 118608 57990
rect 51998 57874 52050 57886
rect 51998 57810 52050 57822
rect 52446 57874 52498 57886
rect 52446 57810 52498 57822
rect 56030 57874 56082 57886
rect 56030 57810 56082 57822
rect 56702 57874 56754 57886
rect 56702 57810 56754 57822
rect 62862 57874 62914 57886
rect 62862 57810 62914 57822
rect 70814 57874 70866 57886
rect 70814 57810 70866 57822
rect 49534 57762 49586 57774
rect 49534 57698 49586 57710
rect 54350 57762 54402 57774
rect 60622 57762 60674 57774
rect 57586 57710 57598 57762
rect 57650 57710 57662 57762
rect 54350 57698 54402 57710
rect 60622 57698 60674 57710
rect 63982 57762 64034 57774
rect 63982 57698 64034 57710
rect 70702 57762 70754 57774
rect 70702 57698 70754 57710
rect 117070 57762 117122 57774
rect 117070 57698 117122 57710
rect 49870 57650 49922 57662
rect 49870 57586 49922 57598
rect 52894 57650 52946 57662
rect 63646 57650 63698 57662
rect 57474 57598 57486 57650
rect 57538 57598 57550 57650
rect 59490 57598 59502 57650
rect 59554 57598 59566 57650
rect 62290 57598 62302 57650
rect 62354 57598 62366 57650
rect 52894 57586 52946 57598
rect 63646 57586 63698 57598
rect 64094 57650 64146 57662
rect 64094 57586 64146 57598
rect 64430 57650 64482 57662
rect 69134 57650 69186 57662
rect 64642 57598 64654 57650
rect 64706 57598 64718 57650
rect 65762 57598 65774 57650
rect 65826 57598 65838 57650
rect 64430 57586 64482 57598
rect 69134 57586 69186 57598
rect 69470 57650 69522 57662
rect 69470 57586 69522 57598
rect 69694 57650 69746 57662
rect 70242 57598 70254 57650
rect 70306 57598 70318 57650
rect 70466 57598 70478 57650
rect 70530 57598 70542 57650
rect 117282 57598 117294 57650
rect 117346 57598 117358 57650
rect 69694 57586 69746 57598
rect 47854 57538 47906 57550
rect 47854 57474 47906 57486
rect 48414 57538 48466 57550
rect 48414 57474 48466 57486
rect 48750 57538 48802 57550
rect 48750 57474 48802 57486
rect 50542 57538 50594 57550
rect 50542 57474 50594 57486
rect 50990 57538 51042 57550
rect 50990 57474 51042 57486
rect 51438 57538 51490 57550
rect 51438 57474 51490 57486
rect 53454 57538 53506 57550
rect 53454 57474 53506 57486
rect 54686 57538 54738 57550
rect 54686 57474 54738 57486
rect 55246 57538 55298 57550
rect 55246 57474 55298 57486
rect 55582 57538 55634 57550
rect 61854 57538 61906 57550
rect 60162 57486 60174 57538
rect 60226 57486 60238 57538
rect 55582 57474 55634 57486
rect 61854 57474 61906 57486
rect 63310 57538 63362 57550
rect 63310 57474 63362 57486
rect 63534 57538 63586 57550
rect 69582 57538 69634 57550
rect 66434 57486 66446 57538
rect 66498 57486 66510 57538
rect 68562 57486 68574 57538
rect 68626 57486 68638 57538
rect 63534 57474 63586 57486
rect 69582 57474 69634 57486
rect 71150 57538 71202 57550
rect 71150 57474 71202 57486
rect 71598 57538 71650 57550
rect 71598 57474 71650 57486
rect 116510 57538 116562 57550
rect 116510 57474 116562 57486
rect 1344 57258 118608 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 96638 57258
rect 96690 57206 96742 57258
rect 96794 57206 96846 57258
rect 96898 57206 118608 57258
rect 1344 57172 118608 57206
rect 65326 57090 65378 57102
rect 41122 57038 41134 57090
rect 41186 57087 41198 57090
rect 41458 57087 41470 57090
rect 41186 57041 41470 57087
rect 41186 57038 41198 57041
rect 41458 57038 41470 57041
rect 41522 57038 41534 57090
rect 65326 57026 65378 57038
rect 41134 56978 41186 56990
rect 58046 56978 58098 56990
rect 56690 56926 56702 56978
rect 56754 56926 56766 56978
rect 41134 56914 41186 56926
rect 58046 56914 58098 56926
rect 58494 56978 58546 56990
rect 58494 56914 58546 56926
rect 58942 56978 58994 56990
rect 58942 56914 58994 56926
rect 59278 56978 59330 56990
rect 59278 56914 59330 56926
rect 59838 56978 59890 56990
rect 59838 56914 59890 56926
rect 59950 56978 60002 56990
rect 59950 56914 60002 56926
rect 61966 56978 62018 56990
rect 61966 56914 62018 56926
rect 62638 56978 62690 56990
rect 62638 56914 62690 56926
rect 64430 56978 64482 56990
rect 66222 56978 66274 56990
rect 69246 56978 69298 56990
rect 65538 56926 65550 56978
rect 65602 56926 65614 56978
rect 66994 56926 67006 56978
rect 67058 56926 67070 56978
rect 70914 56926 70926 56978
rect 70978 56926 70990 56978
rect 73042 56926 73054 56978
rect 73106 56926 73118 56978
rect 64430 56914 64482 56926
rect 66222 56914 66274 56926
rect 69246 56914 69298 56926
rect 41694 56866 41746 56878
rect 47406 56866 47458 56878
rect 52670 56866 52722 56878
rect 57262 56866 57314 56878
rect 3042 56814 3054 56866
rect 3106 56814 3118 56866
rect 45938 56814 45950 56866
rect 46002 56814 46014 56866
rect 48514 56814 48526 56866
rect 48578 56814 48590 56866
rect 53890 56814 53902 56866
rect 53954 56814 53966 56866
rect 41694 56802 41746 56814
rect 47406 56802 47458 56814
rect 52670 56802 52722 56814
rect 57262 56802 57314 56814
rect 57598 56866 57650 56878
rect 64318 56866 64370 56878
rect 63970 56814 63982 56866
rect 64034 56814 64046 56866
rect 57598 56802 57650 56814
rect 64318 56802 64370 56814
rect 67902 56866 67954 56878
rect 70242 56814 70254 56866
rect 70306 56814 70318 56866
rect 67902 56802 67954 56814
rect 42254 56754 42306 56766
rect 66670 56754 66722 56766
rect 1922 56702 1934 56754
rect 1986 56702 1998 56754
rect 49186 56702 49198 56754
rect 49250 56702 49262 56754
rect 54562 56702 54574 56754
rect 54626 56702 54638 56754
rect 42254 56690 42306 56702
rect 66670 56690 66722 56702
rect 3502 56642 3554 56654
rect 3502 56578 3554 56590
rect 46174 56642 46226 56654
rect 46174 56578 46226 56590
rect 46958 56642 47010 56654
rect 46958 56578 47010 56590
rect 47966 56642 48018 56654
rect 52222 56642 52274 56654
rect 51426 56590 51438 56642
rect 51490 56590 51502 56642
rect 47966 56578 48018 56590
rect 52222 56578 52274 56590
rect 57374 56642 57426 56654
rect 57374 56578 57426 56590
rect 60062 56642 60114 56654
rect 60062 56578 60114 56590
rect 60734 56642 60786 56654
rect 60734 56578 60786 56590
rect 61518 56642 61570 56654
rect 61518 56578 61570 56590
rect 65550 56642 65602 56654
rect 65550 56578 65602 56590
rect 66894 56642 66946 56654
rect 66894 56578 66946 56590
rect 67454 56642 67506 56654
rect 67454 56578 67506 56590
rect 68574 56642 68626 56654
rect 68574 56578 68626 56590
rect 73502 56642 73554 56654
rect 73502 56578 73554 56590
rect 118078 56642 118130 56654
rect 118078 56578 118130 56590
rect 1344 56474 118608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 111998 56474
rect 112050 56422 112102 56474
rect 112154 56422 112206 56474
rect 112258 56422 118608 56474
rect 1344 56388 118608 56422
rect 50094 56306 50146 56318
rect 50094 56242 50146 56254
rect 53790 56306 53842 56318
rect 57934 56306 57986 56318
rect 55010 56254 55022 56306
rect 55074 56254 55086 56306
rect 53790 56242 53842 56254
rect 57934 56242 57986 56254
rect 58606 56306 58658 56318
rect 58606 56242 58658 56254
rect 60174 56306 60226 56318
rect 60174 56242 60226 56254
rect 62414 56306 62466 56318
rect 62414 56242 62466 56254
rect 64318 56306 64370 56318
rect 64318 56242 64370 56254
rect 65438 56306 65490 56318
rect 65438 56242 65490 56254
rect 67790 56306 67842 56318
rect 67790 56242 67842 56254
rect 68462 56306 68514 56318
rect 68462 56242 68514 56254
rect 68574 56306 68626 56318
rect 68574 56242 68626 56254
rect 68686 56306 68738 56318
rect 68686 56242 68738 56254
rect 49646 56194 49698 56206
rect 47058 56142 47070 56194
rect 47122 56142 47134 56194
rect 49646 56130 49698 56142
rect 51102 56194 51154 56206
rect 51102 56130 51154 56142
rect 54462 56194 54514 56206
rect 54462 56130 54514 56142
rect 55358 56194 55410 56206
rect 55358 56130 55410 56142
rect 56142 56194 56194 56206
rect 56142 56130 56194 56142
rect 59054 56194 59106 56206
rect 59054 56130 59106 56142
rect 59726 56194 59778 56206
rect 59726 56130 59778 56142
rect 63534 56194 63586 56206
rect 63534 56130 63586 56142
rect 63758 56194 63810 56206
rect 63758 56130 63810 56142
rect 80334 56194 80386 56206
rect 80334 56130 80386 56142
rect 114494 56194 114546 56206
rect 114494 56130 114546 56142
rect 48862 56082 48914 56094
rect 47842 56030 47854 56082
rect 47906 56030 47918 56082
rect 48862 56018 48914 56030
rect 50206 56082 50258 56094
rect 52334 56082 52386 56094
rect 50530 56030 50542 56082
rect 50594 56030 50606 56082
rect 50206 56018 50258 56030
rect 52334 56018 52386 56030
rect 54910 56082 54962 56094
rect 55918 56082 55970 56094
rect 55122 56030 55134 56082
rect 55186 56030 55198 56082
rect 54910 56018 54962 56030
rect 55918 56018 55970 56030
rect 56478 56082 56530 56094
rect 56478 56018 56530 56030
rect 57598 56082 57650 56094
rect 57598 56018 57650 56030
rect 59278 56082 59330 56094
rect 59278 56018 59330 56030
rect 59502 56082 59554 56094
rect 59502 56018 59554 56030
rect 60846 56082 60898 56094
rect 66558 56082 66610 56094
rect 61282 56030 61294 56082
rect 61346 56030 61358 56082
rect 60846 56018 60898 56030
rect 66558 56018 66610 56030
rect 66670 56082 66722 56094
rect 66670 56018 66722 56030
rect 66782 56082 66834 56094
rect 66782 56018 66834 56030
rect 67118 56082 67170 56094
rect 67118 56018 67170 56030
rect 68350 56082 68402 56094
rect 79438 56082 79490 56094
rect 68898 56030 68910 56082
rect 68962 56030 68974 56082
rect 70130 56030 70142 56082
rect 70194 56030 70206 56082
rect 68350 56018 68402 56030
rect 79438 56018 79490 56030
rect 79998 56082 80050 56094
rect 114930 56030 114942 56082
rect 114994 56030 115006 56082
rect 79998 56018 80050 56030
rect 48302 55970 48354 55982
rect 44930 55918 44942 55970
rect 44994 55918 45006 55970
rect 48302 55906 48354 55918
rect 49870 55970 49922 55982
rect 49870 55906 49922 55918
rect 51438 55970 51490 55982
rect 51438 55906 51490 55918
rect 51886 55970 51938 55982
rect 51886 55906 51938 55918
rect 52894 55970 52946 55982
rect 52894 55906 52946 55918
rect 53678 55970 53730 55982
rect 53678 55906 53730 55918
rect 54686 55970 54738 55982
rect 54686 55906 54738 55918
rect 56366 55970 56418 55982
rect 56366 55906 56418 55918
rect 61742 55970 61794 55982
rect 61742 55906 61794 55918
rect 62862 55970 62914 55982
rect 62862 55906 62914 55918
rect 63646 55970 63698 55982
rect 63646 55906 63698 55918
rect 65774 55970 65826 55982
rect 65774 55906 65826 55918
rect 67342 55970 67394 55982
rect 67342 55906 67394 55918
rect 67790 55970 67842 55982
rect 67790 55906 67842 55918
rect 69582 55970 69634 55982
rect 71038 55970 71090 55982
rect 70354 55918 70366 55970
rect 70418 55918 70430 55970
rect 69582 55906 69634 55918
rect 71038 55906 71090 55918
rect 71486 55970 71538 55982
rect 71486 55906 71538 55918
rect 71934 55970 71986 55982
rect 115826 55918 115838 55970
rect 115890 55918 115902 55970
rect 71934 55906 71986 55918
rect 50094 55858 50146 55870
rect 53454 55858 53506 55870
rect 50754 55806 50766 55858
rect 50818 55855 50830 55858
rect 51874 55855 51886 55858
rect 50818 55809 51886 55855
rect 50818 55806 50830 55809
rect 51874 55806 51886 55809
rect 51938 55855 51950 55858
rect 53106 55855 53118 55858
rect 51938 55809 53118 55855
rect 51938 55806 51950 55809
rect 53106 55806 53118 55809
rect 53170 55806 53182 55858
rect 50094 55794 50146 55806
rect 53454 55794 53506 55806
rect 53790 55858 53842 55870
rect 53790 55794 53842 55806
rect 59166 55858 59218 55870
rect 59166 55794 59218 55806
rect 1344 55690 118608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 118608 55690
rect 1344 55604 118608 55638
rect 40910 55522 40962 55534
rect 40910 55458 40962 55470
rect 46398 55522 46450 55534
rect 46398 55458 46450 55470
rect 49646 55522 49698 55534
rect 49646 55458 49698 55470
rect 49982 55522 50034 55534
rect 49982 55458 50034 55470
rect 55022 55522 55074 55534
rect 67778 55470 67790 55522
rect 67842 55519 67854 55522
rect 68226 55519 68238 55522
rect 67842 55473 68238 55519
rect 67842 55470 67854 55473
rect 68226 55470 68238 55473
rect 68290 55470 68302 55522
rect 55022 55458 55074 55470
rect 40014 55410 40066 55422
rect 40014 55346 40066 55358
rect 52558 55410 52610 55422
rect 52558 55346 52610 55358
rect 54126 55410 54178 55422
rect 54126 55346 54178 55358
rect 56814 55410 56866 55422
rect 56814 55346 56866 55358
rect 57486 55410 57538 55422
rect 57486 55346 57538 55358
rect 58942 55410 58994 55422
rect 58942 55346 58994 55358
rect 59390 55410 59442 55422
rect 59390 55346 59442 55358
rect 60062 55410 60114 55422
rect 60062 55346 60114 55358
rect 61294 55410 61346 55422
rect 61294 55346 61346 55358
rect 62078 55410 62130 55422
rect 62078 55346 62130 55358
rect 64206 55410 64258 55422
rect 64206 55346 64258 55358
rect 64654 55410 64706 55422
rect 64654 55346 64706 55358
rect 65550 55410 65602 55422
rect 65550 55346 65602 55358
rect 65998 55410 66050 55422
rect 65998 55346 66050 55358
rect 67342 55410 67394 55422
rect 67342 55346 67394 55358
rect 67790 55410 67842 55422
rect 67790 55346 67842 55358
rect 68574 55410 68626 55422
rect 115826 55358 115838 55410
rect 115890 55358 115902 55410
rect 68574 55346 68626 55358
rect 40798 55298 40850 55310
rect 40798 55234 40850 55246
rect 46734 55298 46786 55310
rect 49198 55298 49250 55310
rect 47506 55246 47518 55298
rect 47570 55246 47582 55298
rect 46734 55234 46786 55246
rect 49198 55234 49250 55246
rect 50542 55298 50594 55310
rect 50542 55234 50594 55246
rect 51214 55298 51266 55310
rect 51214 55234 51266 55246
rect 51550 55298 51602 55310
rect 51550 55234 51602 55246
rect 52334 55298 52386 55310
rect 52334 55234 52386 55246
rect 52782 55298 52834 55310
rect 52782 55234 52834 55246
rect 53678 55298 53730 55310
rect 53678 55234 53730 55246
rect 53902 55298 53954 55310
rect 55134 55298 55186 55310
rect 59166 55298 59218 55310
rect 54674 55246 54686 55298
rect 54738 55295 54750 55298
rect 54898 55295 54910 55298
rect 54738 55249 54910 55295
rect 54738 55246 54750 55249
rect 54898 55246 54910 55249
rect 54962 55246 54974 55298
rect 57922 55246 57934 55298
rect 57986 55246 57998 55298
rect 53902 55234 53954 55246
rect 55134 55234 55186 55246
rect 59166 55234 59218 55246
rect 59502 55298 59554 55310
rect 59502 55234 59554 55246
rect 61854 55298 61906 55310
rect 62526 55298 62578 55310
rect 62290 55246 62302 55298
rect 62354 55246 62366 55298
rect 61854 55234 61906 55246
rect 62526 55234 62578 55246
rect 62862 55298 62914 55310
rect 62862 55234 62914 55246
rect 68238 55298 68290 55310
rect 68238 55234 68290 55246
rect 69694 55298 69746 55310
rect 69694 55234 69746 55246
rect 70030 55298 70082 55310
rect 70030 55234 70082 55246
rect 70366 55298 70418 55310
rect 70366 55234 70418 55246
rect 70590 55298 70642 55310
rect 70590 55234 70642 55246
rect 71486 55298 71538 55310
rect 114930 55246 114942 55298
rect 114994 55246 115006 55298
rect 71486 55234 71538 55246
rect 50990 55186 51042 55198
rect 47282 55134 47294 55186
rect 47346 55134 47358 55186
rect 50990 55122 51042 55134
rect 52110 55186 52162 55198
rect 52110 55122 52162 55134
rect 53454 55186 53506 55198
rect 53454 55122 53506 55134
rect 58270 55186 58322 55198
rect 58270 55122 58322 55134
rect 62974 55186 63026 55198
rect 62974 55122 63026 55134
rect 69582 55186 69634 55198
rect 69582 55122 69634 55134
rect 71038 55186 71090 55198
rect 71038 55122 71090 55134
rect 1822 55074 1874 55086
rect 1822 55010 1874 55022
rect 39678 55074 39730 55086
rect 39678 55010 39730 55022
rect 40686 55074 40738 55086
rect 40686 55010 40738 55022
rect 45838 55074 45890 55086
rect 45838 55010 45890 55022
rect 48190 55074 48242 55086
rect 48190 55010 48242 55022
rect 48638 55074 48690 55086
rect 48638 55010 48690 55022
rect 49758 55074 49810 55086
rect 49758 55010 49810 55022
rect 51438 55074 51490 55086
rect 51438 55010 51490 55022
rect 54574 55074 54626 55086
rect 54574 55010 54626 55022
rect 55246 55074 55298 55086
rect 55246 55010 55298 55022
rect 55918 55074 55970 55086
rect 55918 55010 55970 55022
rect 56254 55074 56306 55086
rect 56254 55010 56306 55022
rect 58158 55074 58210 55086
rect 58158 55010 58210 55022
rect 59054 55074 59106 55086
rect 59054 55010 59106 55022
rect 60622 55074 60674 55086
rect 60622 55010 60674 55022
rect 62302 55074 62354 55086
rect 62302 55010 62354 55022
rect 63534 55074 63586 55086
rect 63534 55010 63586 55022
rect 65102 55074 65154 55086
rect 65102 55010 65154 55022
rect 66446 55074 66498 55086
rect 66446 55010 66498 55022
rect 69470 55074 69522 55086
rect 69470 55010 69522 55022
rect 70366 55074 70418 55086
rect 70366 55010 70418 55022
rect 71934 55074 71986 55086
rect 71934 55010 71986 55022
rect 114382 55074 114434 55086
rect 114382 55010 114434 55022
rect 1344 54906 118608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 111998 54906
rect 112050 54854 112102 54906
rect 112154 54854 112206 54906
rect 112258 54854 118608 54906
rect 1344 54820 118608 54854
rect 40798 54738 40850 54750
rect 40798 54674 40850 54686
rect 41694 54738 41746 54750
rect 41694 54674 41746 54686
rect 45726 54738 45778 54750
rect 45726 54674 45778 54686
rect 46510 54738 46562 54750
rect 46510 54674 46562 54686
rect 47854 54738 47906 54750
rect 47854 54674 47906 54686
rect 48862 54738 48914 54750
rect 48862 54674 48914 54686
rect 51886 54738 51938 54750
rect 51886 54674 51938 54686
rect 53006 54738 53058 54750
rect 53006 54674 53058 54686
rect 53902 54738 53954 54750
rect 53902 54674 53954 54686
rect 56702 54738 56754 54750
rect 56702 54674 56754 54686
rect 59166 54738 59218 54750
rect 59166 54674 59218 54686
rect 64430 54738 64482 54750
rect 64430 54674 64482 54686
rect 68686 54738 68738 54750
rect 68686 54674 68738 54686
rect 41582 54626 41634 54638
rect 41582 54562 41634 54574
rect 41806 54626 41858 54638
rect 41806 54562 41858 54574
rect 46174 54626 46226 54638
rect 46174 54562 46226 54574
rect 49534 54626 49586 54638
rect 63646 54626 63698 54638
rect 51426 54574 51438 54626
rect 51490 54623 51502 54626
rect 51762 54623 51774 54626
rect 51490 54577 51774 54623
rect 51490 54574 51502 54577
rect 51762 54574 51774 54577
rect 51826 54574 51838 54626
rect 49534 54562 49586 54574
rect 63646 54562 63698 54574
rect 63870 54626 63922 54638
rect 63870 54562 63922 54574
rect 66558 54626 66610 54638
rect 66558 54562 66610 54574
rect 67902 54626 67954 54638
rect 67902 54562 67954 54574
rect 68126 54626 68178 54638
rect 68126 54562 68178 54574
rect 89966 54626 90018 54638
rect 89966 54562 90018 54574
rect 47406 54514 47458 54526
rect 47406 54450 47458 54462
rect 49870 54514 49922 54526
rect 49870 54450 49922 54462
rect 50206 54514 50258 54526
rect 50206 54450 50258 54462
rect 51214 54514 51266 54526
rect 52222 54514 52274 54526
rect 51762 54462 51774 54514
rect 51826 54462 51838 54514
rect 51214 54450 51266 54462
rect 52222 54450 52274 54462
rect 54574 54514 54626 54526
rect 54574 54450 54626 54462
rect 55022 54514 55074 54526
rect 55022 54450 55074 54462
rect 57598 54514 57650 54526
rect 58494 54514 58546 54526
rect 89630 54514 89682 54526
rect 57810 54462 57822 54514
rect 57874 54462 57886 54514
rect 59378 54462 59390 54514
rect 59442 54462 59454 54514
rect 59938 54462 59950 54514
rect 60002 54462 60014 54514
rect 69794 54462 69806 54514
rect 69858 54462 69870 54514
rect 57598 54450 57650 54462
rect 58494 54450 58546 54462
rect 89630 54450 89682 54462
rect 40350 54402 40402 54414
rect 40350 54338 40402 54350
rect 47070 54402 47122 54414
rect 47070 54338 47122 54350
rect 48414 54402 48466 54414
rect 48414 54338 48466 54350
rect 49982 54402 50034 54414
rect 49982 54338 50034 54350
rect 50878 54402 50930 54414
rect 50878 54338 50930 54350
rect 52894 54402 52946 54414
rect 52894 54338 52946 54350
rect 54350 54402 54402 54414
rect 54350 54338 54402 54350
rect 55806 54402 55858 54414
rect 55806 54338 55858 54350
rect 56254 54402 56306 54414
rect 65438 54402 65490 54414
rect 60722 54350 60734 54402
rect 60786 54350 60798 54402
rect 62962 54350 62974 54402
rect 63026 54350 63038 54402
rect 56254 54338 56306 54350
rect 65438 54338 65490 54350
rect 67342 54402 67394 54414
rect 67342 54338 67394 54350
rect 69134 54402 69186 54414
rect 73278 54402 73330 54414
rect 70466 54350 70478 54402
rect 70530 54350 70542 54402
rect 72594 54350 72606 54402
rect 72658 54350 72670 54402
rect 69134 54338 69186 54350
rect 73278 54338 73330 54350
rect 88510 54402 88562 54414
rect 88510 54338 88562 54350
rect 51998 54290 52050 54302
rect 45826 54238 45838 54290
rect 45890 54287 45902 54290
rect 46610 54287 46622 54290
rect 45890 54241 46622 54287
rect 45890 54238 45902 54241
rect 46610 54238 46622 54241
rect 46674 54238 46686 54290
rect 51998 54226 52050 54238
rect 54798 54290 54850 54302
rect 54798 54226 54850 54238
rect 55470 54290 55522 54302
rect 59054 54290 59106 54302
rect 56130 54238 56142 54290
rect 56194 54287 56206 54290
rect 56914 54287 56926 54290
rect 56194 54241 56926 54287
rect 56194 54238 56206 54241
rect 56914 54238 56926 54241
rect 56978 54238 56990 54290
rect 55470 54226 55522 54238
rect 59054 54226 59106 54238
rect 63982 54290 64034 54302
rect 63982 54226 64034 54238
rect 68238 54290 68290 54302
rect 68238 54226 68290 54238
rect 1344 54122 118608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 118608 54122
rect 1344 54036 118608 54070
rect 49646 53954 49698 53966
rect 49646 53890 49698 53902
rect 59614 53954 59666 53966
rect 66894 53954 66946 53966
rect 61282 53902 61294 53954
rect 61346 53951 61358 53954
rect 61842 53951 61854 53954
rect 61346 53905 61854 53951
rect 61346 53902 61358 53905
rect 61842 53902 61854 53905
rect 61906 53902 61918 53954
rect 59614 53890 59666 53902
rect 66894 53890 66946 53902
rect 67006 53954 67058 53966
rect 67006 53890 67058 53902
rect 70366 53954 70418 53966
rect 70366 53890 70418 53902
rect 46846 53842 46898 53854
rect 46846 53778 46898 53790
rect 48750 53842 48802 53854
rect 59278 53842 59330 53854
rect 68126 53842 68178 53854
rect 54002 53790 54014 53842
rect 54066 53790 54078 53842
rect 63970 53790 63982 53842
rect 64034 53790 64046 53842
rect 70130 53790 70142 53842
rect 70194 53790 70206 53842
rect 48750 53778 48802 53790
rect 59278 53778 59330 53790
rect 68126 53778 68178 53790
rect 45950 53730 46002 53742
rect 49422 53730 49474 53742
rect 48402 53678 48414 53730
rect 48466 53678 48478 53730
rect 45950 53666 46002 53678
rect 49422 53666 49474 53678
rect 49758 53730 49810 53742
rect 49758 53666 49810 53678
rect 50206 53730 50258 53742
rect 50206 53666 50258 53678
rect 50990 53730 51042 53742
rect 50990 53666 51042 53678
rect 51886 53730 51938 53742
rect 60510 53730 60562 53742
rect 58706 53678 58718 53730
rect 58770 53678 58782 53730
rect 51886 53666 51938 53678
rect 60510 53666 60562 53678
rect 61742 53730 61794 53742
rect 61742 53666 61794 53678
rect 62638 53730 62690 53742
rect 67230 53730 67282 53742
rect 63298 53678 63310 53730
rect 63362 53678 63374 53730
rect 62638 53666 62690 53678
rect 67230 53666 67282 53678
rect 67342 53730 67394 53742
rect 71262 53730 71314 53742
rect 70018 53678 70030 53730
rect 70082 53678 70094 53730
rect 67342 53666 67394 53678
rect 71262 53666 71314 53678
rect 45390 53618 45442 53630
rect 45390 53554 45442 53566
rect 48190 53618 48242 53630
rect 48190 53554 48242 53566
rect 48638 53618 48690 53630
rect 48638 53554 48690 53566
rect 49198 53618 49250 53630
rect 49198 53554 49250 53566
rect 50542 53618 50594 53630
rect 50542 53554 50594 53566
rect 51662 53618 51714 53630
rect 51662 53554 51714 53566
rect 51774 53618 51826 53630
rect 51774 53554 51826 53566
rect 62190 53618 62242 53630
rect 62190 53554 62242 53566
rect 68014 53618 68066 53630
rect 68014 53554 68066 53566
rect 46398 53506 46450 53518
rect 46398 53442 46450 53454
rect 47294 53506 47346 53518
rect 47294 53442 47346 53454
rect 47630 53506 47682 53518
rect 47630 53442 47682 53454
rect 49646 53506 49698 53518
rect 59502 53506 59554 53518
rect 52322 53454 52334 53506
rect 52386 53454 52398 53506
rect 49646 53442 49698 53454
rect 59502 53442 59554 53454
rect 60062 53506 60114 53518
rect 60062 53442 60114 53454
rect 61294 53506 61346 53518
rect 68238 53506 68290 53518
rect 66210 53454 66222 53506
rect 66274 53454 66286 53506
rect 61294 53442 61346 53454
rect 68238 53442 68290 53454
rect 69246 53506 69298 53518
rect 69246 53442 69298 53454
rect 70926 53506 70978 53518
rect 70926 53442 70978 53454
rect 1344 53338 118608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 111998 53338
rect 112050 53286 112102 53338
rect 112154 53286 112206 53338
rect 112258 53286 118608 53338
rect 1344 53252 118608 53286
rect 33966 53170 34018 53182
rect 33966 53106 34018 53118
rect 42478 53170 42530 53182
rect 51326 53170 51378 53182
rect 45714 53118 45726 53170
rect 45778 53118 45790 53170
rect 42478 53106 42530 53118
rect 51326 53106 51378 53118
rect 54686 53170 54738 53182
rect 54686 53106 54738 53118
rect 55582 53170 55634 53182
rect 55582 53106 55634 53118
rect 57934 53170 57986 53182
rect 57934 53106 57986 53118
rect 58494 53170 58546 53182
rect 58494 53106 58546 53118
rect 59390 53170 59442 53182
rect 59390 53106 59442 53118
rect 61854 53170 61906 53182
rect 61854 53106 61906 53118
rect 66222 53170 66274 53182
rect 66222 53106 66274 53118
rect 43150 53058 43202 53070
rect 43150 52994 43202 53006
rect 43374 53058 43426 53070
rect 43374 52994 43426 53006
rect 51886 53058 51938 53070
rect 58046 53058 58098 53070
rect 54002 53006 54014 53058
rect 54066 53006 54078 53058
rect 51886 52994 51938 53006
rect 58046 52994 58098 53006
rect 60510 53058 60562 53070
rect 68562 53006 68574 53058
rect 68626 53006 68638 53058
rect 116274 53006 116286 53058
rect 116338 53006 116350 53058
rect 60510 52994 60562 53006
rect 49758 52946 49810 52958
rect 53678 52946 53730 52958
rect 33730 52894 33742 52946
rect 33794 52894 33806 52946
rect 48738 52894 48750 52946
rect 48802 52894 48814 52946
rect 50418 52894 50430 52946
rect 50482 52894 50494 52946
rect 49758 52882 49810 52894
rect 53678 52882 53730 52894
rect 56030 52946 56082 52958
rect 56030 52882 56082 52894
rect 56254 52946 56306 52958
rect 56254 52882 56306 52894
rect 56702 52946 56754 52958
rect 56702 52882 56754 52894
rect 58158 52946 58210 52958
rect 61406 52946 61458 52958
rect 58706 52894 58718 52946
rect 58770 52894 58782 52946
rect 58158 52882 58210 52894
rect 61406 52882 61458 52894
rect 63870 52946 63922 52958
rect 63870 52882 63922 52894
rect 65774 52946 65826 52958
rect 65774 52882 65826 52894
rect 66334 52946 66386 52958
rect 66334 52882 66386 52894
rect 66446 52946 66498 52958
rect 67778 52894 67790 52946
rect 67842 52894 67854 52946
rect 66446 52882 66498 52894
rect 34414 52834 34466 52846
rect 34414 52770 34466 52782
rect 42030 52834 42082 52846
rect 42030 52770 42082 52782
rect 43262 52834 43314 52846
rect 52334 52834 52386 52846
rect 47954 52782 47966 52834
rect 48018 52782 48030 52834
rect 43262 52770 43314 52782
rect 52334 52770 52386 52782
rect 52782 52834 52834 52846
rect 52782 52770 52834 52782
rect 53230 52834 53282 52846
rect 53230 52770 53282 52782
rect 54798 52834 54850 52846
rect 54798 52770 54850 52782
rect 57374 52834 57426 52846
rect 57374 52770 57426 52782
rect 57710 52834 57762 52846
rect 60062 52834 60114 52846
rect 59266 52782 59278 52834
rect 59330 52782 59342 52834
rect 57710 52770 57762 52782
rect 60062 52770 60114 52782
rect 60958 52834 61010 52846
rect 60958 52770 61010 52782
rect 62302 52834 62354 52846
rect 62302 52770 62354 52782
rect 63310 52834 63362 52846
rect 63310 52770 63362 52782
rect 64542 52834 64594 52846
rect 64542 52770 64594 52782
rect 65326 52834 65378 52846
rect 66894 52834 66946 52846
rect 65538 52782 65550 52834
rect 65602 52831 65614 52834
rect 65762 52831 65774 52834
rect 65602 52785 65774 52831
rect 65602 52782 65614 52785
rect 65762 52782 65774 52785
rect 65826 52782 65838 52834
rect 65326 52770 65378 52782
rect 66894 52770 66946 52782
rect 70702 52834 70754 52846
rect 116846 52834 116898 52846
rect 114930 52782 114942 52834
rect 114994 52782 115006 52834
rect 70702 52770 70754 52782
rect 116846 52770 116898 52782
rect 54910 52722 54962 52734
rect 49858 52670 49870 52722
rect 49922 52670 49934 52722
rect 52322 52670 52334 52722
rect 52386 52719 52398 52722
rect 53330 52719 53342 52722
rect 52386 52673 53342 52719
rect 52386 52670 52398 52673
rect 53330 52670 53342 52673
rect 53394 52670 53406 52722
rect 54910 52658 54962 52670
rect 56478 52722 56530 52734
rect 56478 52658 56530 52670
rect 59614 52722 59666 52734
rect 60722 52670 60734 52722
rect 60786 52719 60798 52722
rect 61394 52719 61406 52722
rect 60786 52673 61406 52719
rect 60786 52670 60798 52673
rect 61394 52670 61406 52673
rect 61458 52670 61470 52722
rect 59614 52658 59666 52670
rect 1344 52554 118608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 118608 52554
rect 1344 52468 118608 52502
rect 49198 52386 49250 52398
rect 46610 52334 46622 52386
rect 46674 52383 46686 52386
rect 48178 52383 48190 52386
rect 46674 52337 48190 52383
rect 46674 52334 46686 52337
rect 48178 52334 48190 52337
rect 48242 52383 48254 52386
rect 48626 52383 48638 52386
rect 48242 52337 48638 52383
rect 48242 52334 48254 52337
rect 48626 52334 48638 52337
rect 48690 52334 48702 52386
rect 49198 52322 49250 52334
rect 49534 52386 49586 52398
rect 49534 52322 49586 52334
rect 50094 52386 50146 52398
rect 50094 52322 50146 52334
rect 50430 52386 50482 52398
rect 50430 52322 50482 52334
rect 52222 52386 52274 52398
rect 52222 52322 52274 52334
rect 55918 52386 55970 52398
rect 55918 52322 55970 52334
rect 56366 52386 56418 52398
rect 56366 52322 56418 52334
rect 60286 52386 60338 52398
rect 60286 52322 60338 52334
rect 60622 52386 60674 52398
rect 60622 52322 60674 52334
rect 62414 52386 62466 52398
rect 62414 52322 62466 52334
rect 67790 52386 67842 52398
rect 67790 52322 67842 52334
rect 46062 52274 46114 52286
rect 3266 52222 3278 52274
rect 3330 52222 3342 52274
rect 46062 52210 46114 52222
rect 47294 52274 47346 52286
rect 47294 52210 47346 52222
rect 47742 52274 47794 52286
rect 47742 52210 47794 52222
rect 48190 52274 48242 52286
rect 48190 52210 48242 52222
rect 51998 52274 52050 52286
rect 51998 52210 52050 52222
rect 56814 52274 56866 52286
rect 56814 52210 56866 52222
rect 57262 52274 57314 52286
rect 57262 52210 57314 52222
rect 57710 52274 57762 52286
rect 57710 52210 57762 52222
rect 58158 52274 58210 52286
rect 58158 52210 58210 52222
rect 63086 52274 63138 52286
rect 63086 52210 63138 52222
rect 64430 52274 64482 52286
rect 64430 52210 64482 52222
rect 65102 52274 65154 52286
rect 65102 52210 65154 52222
rect 67230 52274 67282 52286
rect 67230 52210 67282 52222
rect 68574 52274 68626 52286
rect 68574 52210 68626 52222
rect 69694 52274 69746 52286
rect 74062 52274 74114 52286
rect 73490 52222 73502 52274
rect 73554 52222 73566 52274
rect 69694 52210 69746 52222
rect 74062 52210 74114 52222
rect 46398 52162 46450 52174
rect 46398 52098 46450 52110
rect 48638 52162 48690 52174
rect 48638 52098 48690 52110
rect 51102 52162 51154 52174
rect 51102 52098 51154 52110
rect 54462 52162 54514 52174
rect 55470 52162 55522 52174
rect 54786 52110 54798 52162
rect 54850 52110 54862 52162
rect 54462 52098 54514 52110
rect 55470 52098 55522 52110
rect 55694 52162 55746 52174
rect 69246 52162 69298 52174
rect 61394 52110 61406 52162
rect 61458 52110 61470 52162
rect 63970 52110 63982 52162
rect 64034 52110 64046 52162
rect 65202 52110 65214 52162
rect 65266 52110 65278 52162
rect 66658 52110 66670 52162
rect 66722 52110 66734 52162
rect 66994 52110 67006 52162
rect 67058 52110 67070 52162
rect 70690 52110 70702 52162
rect 70754 52110 70766 52162
rect 55694 52098 55746 52110
rect 69246 52098 69298 52110
rect 54238 52050 54290 52062
rect 1922 51998 1934 52050
rect 1986 51998 1998 52050
rect 54238 51986 54290 51998
rect 59390 52050 59442 52062
rect 59390 51986 59442 51998
rect 64990 52050 65042 52062
rect 64990 51986 65042 51998
rect 65438 52050 65490 52062
rect 71362 51998 71374 52050
rect 71426 51998 71438 52050
rect 65438 51986 65490 51998
rect 46958 51938 47010 51950
rect 46958 51874 47010 51886
rect 49310 51938 49362 51950
rect 49310 51874 49362 51886
rect 50318 51938 50370 51950
rect 50318 51874 50370 51886
rect 50990 51938 51042 51950
rect 53790 51938 53842 51950
rect 52546 51886 52558 51938
rect 52610 51886 52622 51938
rect 50990 51874 51042 51886
rect 53790 51874 53842 51886
rect 58830 51938 58882 51950
rect 58830 51874 58882 51886
rect 58942 51938 58994 51950
rect 58942 51874 58994 51886
rect 59054 51938 59106 51950
rect 59054 51874 59106 51886
rect 59166 51938 59218 51950
rect 59166 51874 59218 51886
rect 60510 51938 60562 51950
rect 60510 51874 60562 51886
rect 67902 51938 67954 51950
rect 67902 51874 67954 51886
rect 68014 51938 68066 51950
rect 68014 51874 68066 51886
rect 1344 51770 118608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 111998 51770
rect 112050 51718 112102 51770
rect 112154 51718 112206 51770
rect 112258 51718 118608 51770
rect 1344 51684 118608 51718
rect 1822 51602 1874 51614
rect 1822 51538 1874 51550
rect 48414 51602 48466 51614
rect 48414 51538 48466 51550
rect 49646 51602 49698 51614
rect 49646 51538 49698 51550
rect 51550 51602 51602 51614
rect 51550 51538 51602 51550
rect 56366 51602 56418 51614
rect 58830 51602 58882 51614
rect 58034 51550 58046 51602
rect 58098 51550 58110 51602
rect 56366 51538 56418 51550
rect 58830 51538 58882 51550
rect 59390 51602 59442 51614
rect 59390 51538 59442 51550
rect 66222 51602 66274 51614
rect 66222 51538 66274 51550
rect 66782 51602 66834 51614
rect 66782 51538 66834 51550
rect 67230 51602 67282 51614
rect 67230 51538 67282 51550
rect 67566 51602 67618 51614
rect 67566 51538 67618 51550
rect 71150 51602 71202 51614
rect 71150 51538 71202 51550
rect 73278 51602 73330 51614
rect 73278 51538 73330 51550
rect 45054 51490 45106 51502
rect 45054 51426 45106 51438
rect 47518 51490 47570 51502
rect 47518 51426 47570 51438
rect 47742 51490 47794 51502
rect 56254 51490 56306 51502
rect 52882 51438 52894 51490
rect 52946 51438 52958 51490
rect 53890 51438 53902 51490
rect 53954 51438 53966 51490
rect 47742 51426 47794 51438
rect 56254 51426 56306 51438
rect 56478 51490 56530 51502
rect 58606 51490 58658 51502
rect 57474 51438 57486 51490
rect 57538 51438 57550 51490
rect 56478 51426 56530 51438
rect 58606 51426 58658 51438
rect 64542 51490 64594 51502
rect 69470 51490 69522 51502
rect 65426 51438 65438 51490
rect 65490 51438 65502 51490
rect 64542 51426 64594 51438
rect 69470 51426 69522 51438
rect 70926 51490 70978 51502
rect 70926 51426 70978 51438
rect 72046 51490 72098 51502
rect 72046 51426 72098 51438
rect 58942 51378 58994 51390
rect 65774 51378 65826 51390
rect 50866 51326 50878 51378
rect 50930 51326 50942 51378
rect 53106 51326 53118 51378
rect 53170 51326 53182 51378
rect 54002 51326 54014 51378
rect 54066 51326 54078 51378
rect 57698 51326 57710 51378
rect 57762 51326 57774 51378
rect 60274 51326 60286 51378
rect 60338 51326 60350 51378
rect 64082 51326 64094 51378
rect 64146 51326 64158 51378
rect 58942 51314 58994 51326
rect 65774 51314 65826 51326
rect 68126 51378 68178 51390
rect 68126 51314 68178 51326
rect 68910 51378 68962 51390
rect 68910 51314 68962 51326
rect 71150 51378 71202 51390
rect 71150 51314 71202 51326
rect 71486 51378 71538 51390
rect 71486 51314 71538 51326
rect 72158 51378 72210 51390
rect 72370 51326 72382 51378
rect 72434 51326 72446 51378
rect 72158 51314 72210 51326
rect 45502 51266 45554 51278
rect 45502 51202 45554 51214
rect 46062 51266 46114 51278
rect 46062 51202 46114 51214
rect 46510 51266 46562 51278
rect 46510 51202 46562 51214
rect 46958 51266 47010 51278
rect 46958 51202 47010 51214
rect 47630 51266 47682 51278
rect 47630 51202 47682 51214
rect 48302 51266 48354 51278
rect 48302 51202 48354 51214
rect 49982 51266 50034 51278
rect 69918 51266 69970 51278
rect 61058 51214 61070 51266
rect 61122 51214 61134 51266
rect 63298 51214 63310 51266
rect 63362 51214 63374 51266
rect 49982 51202 50034 51214
rect 69918 51202 69970 51214
rect 70478 51266 70530 51278
rect 70478 51202 70530 51214
rect 73726 51266 73778 51278
rect 73726 51202 73778 51214
rect 50542 51154 50594 51166
rect 45602 51102 45614 51154
rect 45666 51151 45678 51154
rect 46498 51151 46510 51154
rect 45666 51105 46510 51151
rect 45666 51102 45678 51105
rect 46498 51102 46510 51105
rect 46562 51102 46574 51154
rect 50542 51090 50594 51102
rect 50878 51154 50930 51166
rect 50878 51090 50930 51102
rect 51438 51154 51490 51166
rect 51438 51090 51490 51102
rect 51774 51154 51826 51166
rect 51774 51090 51826 51102
rect 52446 51154 52498 51166
rect 52446 51090 52498 51102
rect 68798 51154 68850 51166
rect 68798 51090 68850 51102
rect 1344 50986 118608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 118608 50986
rect 1344 50900 118608 50934
rect 54238 50818 54290 50830
rect 53330 50766 53342 50818
rect 53394 50815 53406 50818
rect 53554 50815 53566 50818
rect 53394 50769 53566 50815
rect 53394 50766 53406 50769
rect 53554 50766 53566 50769
rect 53618 50766 53630 50818
rect 61506 50766 61518 50818
rect 61570 50766 61582 50818
rect 67330 50766 67342 50818
rect 67394 50815 67406 50818
rect 68786 50815 68798 50818
rect 67394 50769 68798 50815
rect 67394 50766 67406 50769
rect 68786 50766 68798 50769
rect 68850 50766 68862 50818
rect 54238 50754 54290 50766
rect 49198 50706 49250 50718
rect 45490 50654 45502 50706
rect 45554 50654 45566 50706
rect 49198 50642 49250 50654
rect 50430 50706 50482 50718
rect 50430 50642 50482 50654
rect 52670 50706 52722 50718
rect 52670 50642 52722 50654
rect 53566 50706 53618 50718
rect 60510 50706 60562 50718
rect 55458 50654 55470 50706
rect 55522 50654 55534 50706
rect 56466 50654 56478 50706
rect 56530 50654 56542 50706
rect 58482 50654 58494 50706
rect 58546 50654 58558 50706
rect 59378 50654 59390 50706
rect 59442 50654 59454 50706
rect 53566 50642 53618 50654
rect 60510 50642 60562 50654
rect 64430 50706 64482 50718
rect 64430 50642 64482 50654
rect 65214 50706 65266 50718
rect 65214 50642 65266 50654
rect 67230 50706 67282 50718
rect 67230 50642 67282 50654
rect 68238 50706 68290 50718
rect 68238 50642 68290 50654
rect 68574 50706 68626 50718
rect 72258 50654 72270 50706
rect 72322 50654 72334 50706
rect 115490 50654 115502 50706
rect 115554 50654 115566 50706
rect 68574 50642 68626 50654
rect 50654 50594 50706 50606
rect 51214 50594 51266 50606
rect 48290 50542 48302 50594
rect 48354 50542 48366 50594
rect 50866 50542 50878 50594
rect 50930 50542 50942 50594
rect 50654 50530 50706 50542
rect 51214 50530 51266 50542
rect 52222 50594 52274 50606
rect 59726 50594 59778 50606
rect 54898 50542 54910 50594
rect 54962 50542 54974 50594
rect 56130 50542 56142 50594
rect 56194 50542 56206 50594
rect 58594 50542 58606 50594
rect 58658 50542 58670 50594
rect 52222 50530 52274 50542
rect 59726 50530 59778 50542
rect 59950 50594 60002 50606
rect 63758 50594 63810 50606
rect 65662 50594 65714 50606
rect 62178 50542 62190 50594
rect 62242 50542 62254 50594
rect 64530 50542 64542 50594
rect 64594 50542 64606 50594
rect 59950 50530 60002 50542
rect 63758 50530 63810 50542
rect 65662 50530 65714 50542
rect 66558 50594 66610 50606
rect 66558 50530 66610 50542
rect 67790 50594 67842 50606
rect 72718 50594 72770 50606
rect 69346 50542 69358 50594
rect 69410 50542 69422 50594
rect 116162 50542 116174 50594
rect 116226 50542 116238 50594
rect 117282 50542 117294 50594
rect 117346 50542 117358 50594
rect 67790 50530 67842 50542
rect 72718 50530 72770 50542
rect 50206 50482 50258 50494
rect 47618 50430 47630 50482
rect 47682 50430 47694 50482
rect 50206 50418 50258 50430
rect 51662 50482 51714 50494
rect 51662 50418 51714 50430
rect 51886 50482 51938 50494
rect 51886 50418 51938 50430
rect 54350 50482 54402 50494
rect 64318 50482 64370 50494
rect 117070 50482 117122 50494
rect 55234 50430 55246 50482
rect 55298 50430 55310 50482
rect 61618 50430 61630 50482
rect 61682 50430 61694 50482
rect 70130 50430 70142 50482
rect 70194 50430 70206 50482
rect 54350 50418 54402 50430
rect 64318 50418 64370 50430
rect 117070 50418 117122 50430
rect 49758 50370 49810 50382
rect 51550 50370 51602 50382
rect 50754 50318 50766 50370
rect 50818 50318 50830 50370
rect 49758 50306 49810 50318
rect 51550 50306 51602 50318
rect 54238 50370 54290 50382
rect 64766 50370 64818 50382
rect 63410 50318 63422 50370
rect 63474 50318 63486 50370
rect 54238 50306 54290 50318
rect 64766 50306 64818 50318
rect 66670 50370 66722 50382
rect 66670 50306 66722 50318
rect 66894 50370 66946 50382
rect 66894 50306 66946 50318
rect 1344 50202 118608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 111998 50202
rect 112050 50150 112102 50202
rect 112154 50150 112206 50202
rect 112258 50150 118608 50202
rect 1344 50116 118608 50150
rect 45838 50034 45890 50046
rect 45838 49970 45890 49982
rect 46398 50034 46450 50046
rect 46398 49970 46450 49982
rect 47070 50034 47122 50046
rect 47070 49970 47122 49982
rect 47966 50034 48018 50046
rect 47966 49970 48018 49982
rect 48750 50034 48802 50046
rect 53230 50034 53282 50046
rect 50418 49982 50430 50034
rect 50482 49982 50494 50034
rect 48750 49970 48802 49982
rect 53230 49970 53282 49982
rect 54574 50034 54626 50046
rect 54574 49970 54626 49982
rect 63198 50034 63250 50046
rect 63198 49970 63250 49982
rect 64430 50034 64482 50046
rect 64430 49970 64482 49982
rect 70030 50034 70082 50046
rect 70030 49970 70082 49982
rect 116846 50034 116898 50046
rect 116846 49970 116898 49982
rect 47406 49922 47458 49934
rect 47406 49858 47458 49870
rect 50878 49922 50930 49934
rect 50878 49858 50930 49870
rect 52110 49922 52162 49934
rect 52110 49858 52162 49870
rect 52334 49922 52386 49934
rect 52334 49858 52386 49870
rect 53678 49922 53730 49934
rect 53678 49858 53730 49870
rect 54350 49922 54402 49934
rect 64206 49922 64258 49934
rect 55010 49870 55022 49922
rect 55074 49870 55086 49922
rect 60610 49870 60622 49922
rect 60674 49870 60686 49922
rect 54350 49858 54402 49870
rect 64206 49858 64258 49870
rect 72046 49922 72098 49934
rect 72046 49858 72098 49870
rect 72270 49922 72322 49934
rect 72270 49858 72322 49870
rect 45502 49810 45554 49822
rect 45502 49746 45554 49758
rect 46734 49810 46786 49822
rect 46734 49746 46786 49758
rect 47070 49810 47122 49822
rect 50430 49810 50482 49822
rect 50194 49758 50206 49810
rect 50258 49758 50270 49810
rect 47070 49746 47122 49758
rect 50430 49746 50482 49758
rect 50542 49810 50594 49822
rect 50542 49746 50594 49758
rect 54238 49810 54290 49822
rect 56814 49810 56866 49822
rect 63982 49810 64034 49822
rect 68126 49810 68178 49822
rect 56354 49758 56366 49810
rect 56418 49758 56430 49810
rect 57810 49758 57822 49810
rect 57874 49758 57886 49810
rect 66770 49758 66782 49810
rect 66834 49758 66846 49810
rect 54238 49746 54290 49758
rect 56814 49746 56866 49758
rect 63982 49746 64034 49758
rect 68126 49746 68178 49758
rect 69806 49810 69858 49822
rect 69806 49746 69858 49758
rect 70030 49810 70082 49822
rect 70030 49746 70082 49758
rect 70366 49810 70418 49822
rect 70366 49746 70418 49758
rect 70926 49810 70978 49822
rect 70926 49746 70978 49758
rect 45054 49698 45106 49710
rect 45054 49634 45106 49646
rect 48414 49698 48466 49710
rect 48414 49634 48466 49646
rect 49534 49698 49586 49710
rect 49534 49634 49586 49646
rect 51550 49698 51602 49710
rect 52782 49698 52834 49710
rect 52098 49646 52110 49698
rect 52162 49646 52174 49698
rect 51550 49634 51602 49646
rect 52782 49634 52834 49646
rect 64094 49698 64146 49710
rect 64094 49634 64146 49646
rect 65326 49698 65378 49710
rect 65326 49634 65378 49646
rect 65774 49698 65826 49710
rect 68574 49698 68626 49710
rect 66882 49646 66894 49698
rect 66946 49646 66958 49698
rect 65774 49634 65826 49646
rect 68574 49634 68626 49646
rect 69022 49698 69074 49710
rect 69022 49634 69074 49646
rect 71486 49698 71538 49710
rect 73278 49698 73330 49710
rect 72258 49646 72270 49698
rect 72322 49646 72334 49698
rect 71486 49634 71538 49646
rect 73278 49634 73330 49646
rect 67218 49534 67230 49586
rect 67282 49534 67294 49586
rect 1344 49418 118608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 118608 49418
rect 1344 49332 118608 49366
rect 51102 49250 51154 49262
rect 70578 49198 70590 49250
rect 70642 49247 70654 49250
rect 70914 49247 70926 49250
rect 70642 49201 70926 49247
rect 70642 49198 70654 49201
rect 70914 49198 70926 49201
rect 70978 49198 70990 49250
rect 51102 49186 51154 49198
rect 46510 49138 46562 49150
rect 46510 49074 46562 49086
rect 46958 49138 47010 49150
rect 46958 49074 47010 49086
rect 47854 49138 47906 49150
rect 47854 49074 47906 49086
rect 48414 49138 48466 49150
rect 48414 49074 48466 49086
rect 48862 49138 48914 49150
rect 48862 49074 48914 49086
rect 50318 49138 50370 49150
rect 50318 49074 50370 49086
rect 52670 49138 52722 49150
rect 52670 49074 52722 49086
rect 53454 49138 53506 49150
rect 53454 49074 53506 49086
rect 54126 49138 54178 49150
rect 61518 49138 61570 49150
rect 58818 49086 58830 49138
rect 58882 49086 58894 49138
rect 54126 49074 54178 49086
rect 61518 49074 61570 49086
rect 62974 49138 63026 49150
rect 68014 49138 68066 49150
rect 64642 49086 64654 49138
rect 64706 49086 64718 49138
rect 62974 49074 63026 49086
rect 68014 49074 68066 49086
rect 68350 49138 68402 49150
rect 68350 49074 68402 49086
rect 69582 49138 69634 49150
rect 69582 49074 69634 49086
rect 70590 49138 70642 49150
rect 70590 49074 70642 49086
rect 71822 49138 71874 49150
rect 115490 49086 115502 49138
rect 115554 49086 115566 49138
rect 71822 49074 71874 49086
rect 49534 49026 49586 49038
rect 49298 48974 49310 49026
rect 49362 48974 49374 49026
rect 49534 48962 49586 48974
rect 49646 49026 49698 49038
rect 49646 48962 49698 48974
rect 49982 49026 50034 49038
rect 49982 48962 50034 48974
rect 50542 49026 50594 49038
rect 55246 49026 55298 49038
rect 53890 48974 53902 49026
rect 53954 48974 53966 49026
rect 50542 48962 50594 48974
rect 55246 48962 55298 48974
rect 56478 49026 56530 49038
rect 56478 48962 56530 48974
rect 57486 49026 57538 49038
rect 57486 48962 57538 48974
rect 57710 49026 57762 49038
rect 61630 49026 61682 49038
rect 59938 48974 59950 49026
rect 60002 48974 60014 49026
rect 57710 48962 57762 48974
rect 61630 48962 61682 48974
rect 62078 49026 62130 49038
rect 62078 48962 62130 48974
rect 62862 49026 62914 49038
rect 62862 48962 62914 48974
rect 63198 49026 63250 49038
rect 63858 48974 63870 49026
rect 63922 48974 63934 49026
rect 116162 48974 116174 49026
rect 116226 48974 116238 49026
rect 63198 48962 63250 48974
rect 46062 48914 46114 48926
rect 46062 48850 46114 48862
rect 52110 48914 52162 48926
rect 52110 48850 52162 48862
rect 54238 48914 54290 48926
rect 54238 48850 54290 48862
rect 55134 48914 55186 48926
rect 55134 48850 55186 48862
rect 55358 48914 55410 48926
rect 61406 48914 61458 48926
rect 60050 48862 60062 48914
rect 60114 48862 60126 48914
rect 55358 48850 55410 48862
rect 61406 48850 61458 48862
rect 63086 48914 63138 48926
rect 63086 48850 63138 48862
rect 1822 48802 1874 48814
rect 1822 48738 1874 48750
rect 45726 48802 45778 48814
rect 45726 48738 45778 48750
rect 47406 48802 47458 48814
rect 47406 48738 47458 48750
rect 50318 48802 50370 48814
rect 50318 48738 50370 48750
rect 51214 48802 51266 48814
rect 51214 48738 51266 48750
rect 51326 48802 51378 48814
rect 51326 48738 51378 48750
rect 51998 48802 52050 48814
rect 56926 48802 56978 48814
rect 62750 48802 62802 48814
rect 67454 48802 67506 48814
rect 55794 48750 55806 48802
rect 55858 48750 55870 48802
rect 58034 48750 58046 48802
rect 58098 48750 58110 48802
rect 66882 48750 66894 48802
rect 66946 48750 66958 48802
rect 51998 48738 52050 48750
rect 56926 48738 56978 48750
rect 62750 48738 62802 48750
rect 67454 48738 67506 48750
rect 71038 48802 71090 48814
rect 71038 48738 71090 48750
rect 116958 48802 117010 48814
rect 116958 48738 117010 48750
rect 1344 48634 118608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 111998 48634
rect 112050 48582 112102 48634
rect 112154 48582 112206 48634
rect 112258 48582 118608 48634
rect 1344 48548 118608 48582
rect 45278 48466 45330 48478
rect 45278 48402 45330 48414
rect 48862 48466 48914 48478
rect 48862 48402 48914 48414
rect 56702 48466 56754 48478
rect 64206 48466 64258 48478
rect 58706 48414 58718 48466
rect 58770 48414 58782 48466
rect 56702 48402 56754 48414
rect 64206 48402 64258 48414
rect 65886 48466 65938 48478
rect 65886 48402 65938 48414
rect 67118 48466 67170 48478
rect 67118 48402 67170 48414
rect 67678 48466 67730 48478
rect 67678 48402 67730 48414
rect 117070 48466 117122 48478
rect 117070 48402 117122 48414
rect 46734 48354 46786 48366
rect 46734 48290 46786 48302
rect 47070 48354 47122 48366
rect 47070 48290 47122 48302
rect 47966 48354 48018 48366
rect 47966 48290 48018 48302
rect 49646 48354 49698 48366
rect 49646 48290 49698 48302
rect 49870 48354 49922 48366
rect 49870 48290 49922 48302
rect 51550 48354 51602 48366
rect 51550 48290 51602 48302
rect 53006 48354 53058 48366
rect 53006 48290 53058 48302
rect 58158 48354 58210 48366
rect 61742 48354 61794 48366
rect 58818 48302 58830 48354
rect 58882 48302 58894 48354
rect 58158 48290 58210 48302
rect 61742 48290 61794 48302
rect 67230 48354 67282 48366
rect 67230 48290 67282 48302
rect 68462 48354 68514 48366
rect 68462 48290 68514 48302
rect 47294 48242 47346 48254
rect 47294 48178 47346 48190
rect 49534 48242 49586 48254
rect 52446 48242 52498 48254
rect 57598 48242 57650 48254
rect 52098 48190 52110 48242
rect 52162 48190 52174 48242
rect 55234 48190 55246 48242
rect 55298 48190 55310 48242
rect 49534 48178 49586 48190
rect 52446 48178 52498 48190
rect 57598 48178 57650 48190
rect 59166 48242 59218 48254
rect 59166 48178 59218 48190
rect 59614 48242 59666 48254
rect 63310 48242 63362 48254
rect 60498 48190 60510 48242
rect 60562 48190 60574 48242
rect 61282 48190 61294 48242
rect 61346 48190 61358 48242
rect 61506 48190 61518 48242
rect 61570 48190 61582 48242
rect 63074 48190 63086 48242
rect 63138 48190 63150 48242
rect 59614 48178 59666 48190
rect 63310 48178 63362 48190
rect 63982 48242 64034 48254
rect 63982 48178 64034 48190
rect 64318 48242 64370 48254
rect 67342 48242 67394 48254
rect 70142 48242 70194 48254
rect 66098 48190 66110 48242
rect 66162 48190 66174 48242
rect 67890 48190 67902 48242
rect 67954 48190 67966 48242
rect 68786 48190 68798 48242
rect 68850 48190 68862 48242
rect 116162 48190 116174 48242
rect 116226 48190 116238 48242
rect 117282 48190 117294 48242
rect 117346 48190 117358 48242
rect 64318 48178 64370 48190
rect 67342 48178 67394 48190
rect 70142 48178 70194 48190
rect 45726 48130 45778 48142
rect 45726 48066 45778 48078
rect 46286 48130 46338 48142
rect 46286 48066 46338 48078
rect 46846 48130 46898 48142
rect 55694 48130 55746 48142
rect 47842 48078 47854 48130
rect 47906 48078 47918 48130
rect 50754 48078 50766 48130
rect 50818 48078 50830 48130
rect 54786 48078 54798 48130
rect 54850 48078 54862 48130
rect 46846 48066 46898 48078
rect 55694 48066 55746 48078
rect 56142 48130 56194 48142
rect 56142 48066 56194 48078
rect 58382 48130 58434 48142
rect 61406 48130 61458 48142
rect 60386 48078 60398 48130
rect 60450 48078 60462 48130
rect 58382 48066 58434 48078
rect 61406 48066 61458 48078
rect 66670 48130 66722 48142
rect 66670 48066 66722 48078
rect 67006 48130 67058 48142
rect 69246 48130 69298 48142
rect 68674 48078 68686 48130
rect 68738 48078 68750 48130
rect 67006 48066 67058 48078
rect 69246 48066 69298 48078
rect 69694 48130 69746 48142
rect 69694 48066 69746 48078
rect 70590 48130 70642 48142
rect 115490 48078 115502 48130
rect 115554 48078 115566 48130
rect 70590 48066 70642 48078
rect 48190 48018 48242 48030
rect 48190 47954 48242 47966
rect 58606 48018 58658 48030
rect 65774 48018 65826 48030
rect 63186 47966 63198 48018
rect 63250 47966 63262 48018
rect 58606 47954 58658 47966
rect 65774 47954 65826 47966
rect 1344 47850 118608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 118608 47850
rect 1344 47764 118608 47798
rect 54014 47682 54066 47694
rect 56030 47682 56082 47694
rect 59614 47682 59666 47694
rect 55010 47630 55022 47682
rect 55074 47679 55086 47682
rect 55346 47679 55358 47682
rect 55074 47633 55358 47679
rect 55074 47630 55086 47633
rect 55346 47630 55358 47633
rect 55410 47630 55422 47682
rect 57362 47630 57374 47682
rect 57426 47679 57438 47682
rect 57698 47679 57710 47682
rect 57426 47633 57710 47679
rect 57426 47630 57438 47633
rect 57698 47630 57710 47633
rect 57762 47630 57774 47682
rect 58258 47630 58270 47682
rect 58322 47630 58334 47682
rect 54014 47618 54066 47630
rect 56030 47618 56082 47630
rect 59614 47618 59666 47630
rect 62190 47682 62242 47694
rect 62190 47618 62242 47630
rect 62974 47682 63026 47694
rect 62974 47618 63026 47630
rect 3278 47570 3330 47582
rect 52670 47570 52722 47582
rect 54574 47570 54626 47582
rect 45490 47518 45502 47570
rect 45554 47518 45566 47570
rect 47618 47518 47630 47570
rect 47682 47518 47694 47570
rect 48962 47518 48974 47570
rect 49026 47518 49038 47570
rect 51090 47518 51102 47570
rect 51154 47518 51166 47570
rect 53778 47518 53790 47570
rect 53842 47518 53854 47570
rect 3278 47506 3330 47518
rect 52670 47506 52722 47518
rect 54574 47506 54626 47518
rect 56254 47570 56306 47582
rect 56254 47506 56306 47518
rect 57710 47570 57762 47582
rect 60398 47570 60450 47582
rect 59938 47518 59950 47570
rect 60002 47518 60014 47570
rect 57710 47506 57762 47518
rect 60398 47506 60450 47518
rect 63086 47570 63138 47582
rect 63086 47506 63138 47518
rect 67678 47570 67730 47582
rect 67678 47506 67730 47518
rect 68350 47570 68402 47582
rect 73726 47570 73778 47582
rect 71138 47518 71150 47570
rect 71202 47518 71214 47570
rect 73266 47518 73278 47570
rect 73330 47518 73342 47570
rect 68350 47506 68402 47518
rect 73726 47506 73778 47518
rect 55918 47458 55970 47470
rect 2594 47406 2606 47458
rect 2658 47406 2670 47458
rect 48402 47406 48414 47458
rect 48466 47406 48478 47458
rect 51762 47406 51774 47458
rect 51826 47406 51838 47458
rect 55570 47406 55582 47458
rect 55634 47406 55646 47458
rect 55918 47394 55970 47406
rect 57374 47458 57426 47470
rect 61294 47458 61346 47470
rect 59042 47406 59054 47458
rect 59106 47406 59118 47458
rect 57374 47394 57426 47406
rect 61294 47394 61346 47406
rect 61630 47458 61682 47470
rect 61630 47394 61682 47406
rect 62302 47458 62354 47470
rect 63298 47406 63310 47458
rect 63362 47406 63374 47458
rect 66994 47406 67006 47458
rect 67058 47406 67070 47458
rect 70354 47406 70366 47458
rect 70418 47406 70430 47458
rect 117282 47406 117294 47458
rect 117346 47406 117358 47458
rect 62302 47394 62354 47406
rect 56478 47346 56530 47358
rect 56478 47282 56530 47294
rect 58718 47346 58770 47358
rect 58718 47282 58770 47294
rect 58830 47346 58882 47358
rect 67566 47346 67618 47358
rect 66210 47294 66222 47346
rect 66274 47294 66286 47346
rect 58830 47282 58882 47294
rect 67566 47282 67618 47294
rect 69246 47346 69298 47358
rect 69246 47282 69298 47294
rect 117070 47346 117122 47358
rect 117070 47282 117122 47294
rect 2830 47234 2882 47246
rect 2830 47170 2882 47182
rect 53790 47234 53842 47246
rect 53790 47170 53842 47182
rect 55022 47234 55074 47246
rect 55022 47170 55074 47182
rect 56030 47234 56082 47246
rect 56030 47170 56082 47182
rect 59838 47234 59890 47246
rect 59838 47170 59890 47182
rect 61518 47234 61570 47246
rect 67790 47234 67842 47246
rect 63970 47182 63982 47234
rect 64034 47182 64046 47234
rect 61518 47170 61570 47182
rect 67790 47170 67842 47182
rect 69806 47234 69858 47246
rect 69806 47170 69858 47182
rect 116286 47234 116338 47246
rect 116286 47170 116338 47182
rect 1344 47066 118608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 111998 47066
rect 112050 47014 112102 47066
rect 112154 47014 112206 47066
rect 112258 47014 118608 47066
rect 1344 46980 118608 47014
rect 46846 46898 46898 46910
rect 46846 46834 46898 46846
rect 47518 46898 47570 46910
rect 47518 46834 47570 46846
rect 48750 46898 48802 46910
rect 48750 46834 48802 46846
rect 54350 46898 54402 46910
rect 54350 46834 54402 46846
rect 56590 46898 56642 46910
rect 56590 46834 56642 46846
rect 57374 46898 57426 46910
rect 57374 46834 57426 46846
rect 58270 46898 58322 46910
rect 58270 46834 58322 46846
rect 64094 46898 64146 46910
rect 64094 46834 64146 46846
rect 65326 46898 65378 46910
rect 65326 46834 65378 46846
rect 65774 46898 65826 46910
rect 65774 46834 65826 46846
rect 66670 46898 66722 46910
rect 66670 46834 66722 46846
rect 47294 46786 47346 46798
rect 47294 46722 47346 46734
rect 55806 46786 55858 46798
rect 55806 46722 55858 46734
rect 56030 46786 56082 46798
rect 62638 46786 62690 46798
rect 59938 46734 59950 46786
rect 60002 46734 60014 46786
rect 56030 46722 56082 46734
rect 62638 46722 62690 46734
rect 63198 46786 63250 46798
rect 63198 46722 63250 46734
rect 66222 46786 66274 46798
rect 118078 46786 118130 46798
rect 68674 46734 68686 46786
rect 68738 46734 68750 46786
rect 66222 46722 66274 46734
rect 118078 46722 118130 46734
rect 47630 46674 47682 46686
rect 2818 46622 2830 46674
rect 2882 46622 2894 46674
rect 47630 46610 47682 46622
rect 47854 46674 47906 46686
rect 47854 46610 47906 46622
rect 49870 46674 49922 46686
rect 62862 46674 62914 46686
rect 50530 46622 50542 46674
rect 50594 46622 50606 46674
rect 59266 46622 59278 46674
rect 59330 46622 59342 46674
rect 49870 46610 49922 46622
rect 62862 46610 62914 46622
rect 62974 46674 63026 46686
rect 62974 46610 63026 46622
rect 63086 46674 63138 46686
rect 63086 46610 63138 46622
rect 63758 46674 63810 46686
rect 63758 46610 63810 46622
rect 64094 46674 64146 46686
rect 64094 46610 64146 46622
rect 64318 46674 64370 46686
rect 68002 46622 68014 46674
rect 68066 46622 68078 46674
rect 64318 46610 64370 46622
rect 48414 46562 48466 46574
rect 1922 46510 1934 46562
rect 1986 46510 1998 46562
rect 48414 46498 48466 46510
rect 49982 46562 50034 46574
rect 54686 46562 54738 46574
rect 51314 46510 51326 46562
rect 51378 46510 51390 46562
rect 53442 46510 53454 46562
rect 53506 46510 53518 46562
rect 49982 46498 50034 46510
rect 54686 46498 54738 46510
rect 55134 46562 55186 46574
rect 55134 46498 55186 46510
rect 58606 46562 58658 46574
rect 67230 46562 67282 46574
rect 62066 46510 62078 46562
rect 62130 46510 62142 46562
rect 58606 46498 58658 46510
rect 67230 46498 67282 46510
rect 70814 46562 70866 46574
rect 70814 46498 70866 46510
rect 55694 46450 55746 46462
rect 55694 46386 55746 46398
rect 1344 46282 118608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 118608 46282
rect 1344 46196 118608 46230
rect 50654 46114 50706 46126
rect 52434 46062 52446 46114
rect 52498 46111 52510 46114
rect 52658 46111 52670 46114
rect 52498 46065 52670 46111
rect 52498 46062 52510 46065
rect 52658 46062 52670 46065
rect 52722 46062 52734 46114
rect 59602 46062 59614 46114
rect 59666 46111 59678 46114
rect 59826 46111 59838 46114
rect 59666 46065 59838 46111
rect 59666 46062 59678 46065
rect 59826 46062 59838 46065
rect 59890 46062 59902 46114
rect 50654 46050 50706 46062
rect 50206 46002 50258 46014
rect 52222 46002 52274 46014
rect 45602 45950 45614 46002
rect 45666 45950 45678 46002
rect 47730 45950 47742 46002
rect 47794 45950 47806 46002
rect 50866 45950 50878 46002
rect 50930 45950 50942 46002
rect 50206 45938 50258 45950
rect 52222 45938 52274 45950
rect 52670 46002 52722 46014
rect 52670 45938 52722 45950
rect 53678 46002 53730 46014
rect 60622 46002 60674 46014
rect 55346 45950 55358 46002
rect 55410 45950 55422 46002
rect 53678 45938 53730 45950
rect 60622 45938 60674 45950
rect 67230 46002 67282 46014
rect 115490 45950 115502 46002
rect 115554 45950 115566 46002
rect 67230 45938 67282 45950
rect 54126 45890 54178 45902
rect 58606 45890 58658 45902
rect 3042 45838 3054 45890
rect 3106 45838 3118 45890
rect 48514 45838 48526 45890
rect 48578 45838 48590 45890
rect 54562 45838 54574 45890
rect 54626 45838 54638 45890
rect 54126 45826 54178 45838
rect 58606 45826 58658 45838
rect 58942 45890 58994 45902
rect 61394 45838 61406 45890
rect 61458 45838 61470 45890
rect 116162 45838 116174 45890
rect 116226 45838 116238 45890
rect 58942 45826 58994 45838
rect 68014 45778 68066 45790
rect 1922 45726 1934 45778
rect 1986 45726 1998 45778
rect 63858 45726 63870 45778
rect 63922 45726 63934 45778
rect 68014 45714 68066 45726
rect 3502 45666 3554 45678
rect 3502 45602 3554 45614
rect 49198 45666 49250 45678
rect 49198 45602 49250 45614
rect 49646 45666 49698 45678
rect 49646 45602 49698 45614
rect 50878 45666 50930 45678
rect 50878 45602 50930 45614
rect 51550 45666 51602 45678
rect 58718 45666 58770 45678
rect 57586 45614 57598 45666
rect 57650 45614 57662 45666
rect 51550 45602 51602 45614
rect 58718 45602 58770 45614
rect 59614 45666 59666 45678
rect 59614 45602 59666 45614
rect 60174 45666 60226 45678
rect 60174 45602 60226 45614
rect 67566 45666 67618 45678
rect 67566 45602 67618 45614
rect 1344 45498 118608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 118608 45498
rect 1344 45412 118608 45446
rect 42926 45330 42978 45342
rect 42926 45266 42978 45278
rect 47742 45330 47794 45342
rect 47742 45266 47794 45278
rect 48638 45330 48690 45342
rect 48638 45266 48690 45278
rect 49422 45330 49474 45342
rect 49422 45266 49474 45278
rect 50990 45330 51042 45342
rect 50990 45266 51042 45278
rect 51438 45330 51490 45342
rect 51438 45266 51490 45278
rect 52446 45330 52498 45342
rect 52446 45266 52498 45278
rect 54910 45330 54962 45342
rect 54910 45266 54962 45278
rect 56366 45330 56418 45342
rect 56366 45266 56418 45278
rect 56814 45330 56866 45342
rect 56814 45266 56866 45278
rect 57486 45330 57538 45342
rect 57486 45266 57538 45278
rect 61630 45330 61682 45342
rect 61630 45266 61682 45278
rect 61966 45330 62018 45342
rect 61966 45266 62018 45278
rect 64206 45330 64258 45342
rect 64206 45266 64258 45278
rect 64542 45330 64594 45342
rect 64542 45266 64594 45278
rect 116510 45330 116562 45342
rect 116510 45266 116562 45278
rect 117070 45330 117122 45342
rect 117070 45266 117122 45278
rect 42142 45218 42194 45230
rect 42142 45154 42194 45166
rect 42478 45218 42530 45230
rect 42478 45154 42530 45166
rect 51998 45218 52050 45230
rect 51998 45154 52050 45166
rect 53678 45218 53730 45230
rect 53678 45154 53730 45166
rect 58830 45218 58882 45230
rect 58830 45154 58882 45166
rect 59502 45218 59554 45230
rect 59502 45154 59554 45166
rect 65774 45218 65826 45230
rect 65774 45154 65826 45166
rect 117406 45218 117458 45230
rect 117406 45154 117458 45166
rect 46958 45106 47010 45118
rect 58270 45106 58322 45118
rect 47506 45054 47518 45106
rect 47570 45054 47582 45106
rect 46958 45042 47010 45054
rect 58270 45042 58322 45054
rect 58494 45106 58546 45118
rect 58494 45042 58546 45054
rect 59278 45106 59330 45118
rect 59278 45042 59330 45054
rect 59614 45106 59666 45118
rect 63410 45054 63422 45106
rect 63474 45054 63486 45106
rect 59614 45042 59666 45054
rect 50542 44994 50594 45006
rect 50542 44930 50594 44942
rect 53230 44994 53282 45006
rect 53230 44930 53282 44942
rect 54126 44994 54178 45006
rect 54126 44930 54178 44942
rect 54462 44994 54514 45006
rect 54462 44930 54514 44942
rect 55358 44994 55410 45006
rect 55358 44930 55410 44942
rect 55918 44994 55970 45006
rect 55918 44930 55970 44942
rect 58382 44994 58434 45006
rect 58382 44930 58434 44942
rect 60062 44994 60114 45006
rect 60062 44930 60114 44942
rect 60510 44994 60562 45006
rect 60510 44930 60562 44942
rect 60958 44994 61010 45006
rect 65326 44994 65378 45006
rect 62738 44942 62750 44994
rect 62802 44942 62814 44994
rect 60958 44930 61010 44942
rect 65326 44930 65378 44942
rect 66446 44994 66498 45006
rect 66446 44930 66498 44942
rect 66894 44994 66946 45006
rect 66894 44930 66946 44942
rect 47854 44882 47906 44894
rect 54226 44830 54238 44882
rect 54290 44879 54302 44882
rect 55010 44879 55022 44882
rect 54290 44833 55022 44879
rect 54290 44830 54302 44833
rect 55010 44830 55022 44833
rect 55074 44830 55086 44882
rect 60610 44830 60622 44882
rect 60674 44879 60686 44882
rect 60946 44879 60958 44882
rect 60674 44833 60958 44879
rect 60674 44830 60686 44833
rect 60946 44830 60958 44833
rect 61010 44879 61022 44882
rect 62066 44879 62078 44882
rect 61010 44833 62078 44879
rect 61010 44830 61022 44833
rect 62066 44830 62078 44833
rect 62130 44830 62142 44882
rect 62962 44830 62974 44882
rect 63026 44830 63038 44882
rect 47854 44818 47906 44830
rect 1344 44714 118608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 118608 44714
rect 1344 44628 118608 44662
rect 52110 44546 52162 44558
rect 49074 44494 49086 44546
rect 49138 44543 49150 44546
rect 50306 44543 50318 44546
rect 49138 44497 50318 44543
rect 49138 44494 49150 44497
rect 50306 44494 50318 44497
rect 50370 44494 50382 44546
rect 52110 44482 52162 44494
rect 61966 44546 62018 44558
rect 61966 44482 62018 44494
rect 49086 44434 49138 44446
rect 49086 44370 49138 44382
rect 50430 44434 50482 44446
rect 55918 44434 55970 44446
rect 54226 44382 54238 44434
rect 54290 44382 54302 44434
rect 50430 44370 50482 44382
rect 55918 44370 55970 44382
rect 56702 44434 56754 44446
rect 56702 44370 56754 44382
rect 57374 44434 57426 44446
rect 67902 44434 67954 44446
rect 59490 44382 59502 44434
rect 59554 44382 59566 44434
rect 65090 44382 65102 44434
rect 65154 44382 65166 44434
rect 57374 44370 57426 44382
rect 67902 44370 67954 44382
rect 49982 44322 50034 44334
rect 49982 44258 50034 44270
rect 51886 44322 51938 44334
rect 51886 44258 51938 44270
rect 55022 44322 55074 44334
rect 61294 44322 61346 44334
rect 66110 44322 66162 44334
rect 60274 44270 60286 44322
rect 60338 44270 60350 44322
rect 62402 44270 62414 44322
rect 62466 44270 62478 44322
rect 65650 44270 65662 44322
rect 65714 44270 65726 44322
rect 55022 44258 55074 44270
rect 61294 44258 61346 44270
rect 66110 44258 66162 44270
rect 66894 44322 66946 44334
rect 66894 44258 66946 44270
rect 67230 44322 67282 44334
rect 67230 44258 67282 44270
rect 51326 44210 51378 44222
rect 51326 44146 51378 44158
rect 53678 44210 53730 44222
rect 53678 44146 53730 44158
rect 53790 44210 53842 44222
rect 54798 44210 54850 44222
rect 53890 44158 53902 44210
rect 53954 44158 53966 44210
rect 53790 44146 53842 44158
rect 54798 44146 54850 44158
rect 55358 44210 55410 44222
rect 67454 44210 67506 44222
rect 62962 44158 62974 44210
rect 63026 44158 63038 44210
rect 64194 44158 64206 44210
rect 64258 44158 64270 44210
rect 55358 44146 55410 44158
rect 67454 44146 67506 44158
rect 48078 44098 48130 44110
rect 48078 44034 48130 44046
rect 49534 44098 49586 44110
rect 49534 44034 49586 44046
rect 50878 44098 50930 44110
rect 53454 44098 53506 44110
rect 52434 44046 52446 44098
rect 52498 44046 52510 44098
rect 50878 44034 50930 44046
rect 53454 44034 53506 44046
rect 55134 44098 55186 44110
rect 55134 44034 55186 44046
rect 61630 44098 61682 44110
rect 61630 44034 61682 44046
rect 61854 44098 61906 44110
rect 61854 44034 61906 44046
rect 67006 44098 67058 44110
rect 67006 44034 67058 44046
rect 67118 44098 67170 44110
rect 67118 44034 67170 44046
rect 68462 44098 68514 44110
rect 68462 44034 68514 44046
rect 1344 43930 118608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 118608 43930
rect 1344 43844 118608 43878
rect 59950 43762 60002 43774
rect 64542 43762 64594 43774
rect 61618 43710 61630 43762
rect 61682 43710 61694 43762
rect 59950 43698 60002 43710
rect 64542 43698 64594 43710
rect 68238 43762 68290 43774
rect 68238 43698 68290 43710
rect 52894 43650 52946 43662
rect 57486 43650 57538 43662
rect 54226 43598 54238 43650
rect 54290 43598 54302 43650
rect 52894 43586 52946 43598
rect 57486 43586 57538 43598
rect 63086 43650 63138 43662
rect 63086 43586 63138 43598
rect 63534 43650 63586 43662
rect 63534 43586 63586 43598
rect 66222 43650 66274 43662
rect 116274 43598 116286 43650
rect 116338 43598 116350 43650
rect 66222 43586 66274 43598
rect 50766 43538 50818 43550
rect 58942 43538 58994 43550
rect 50418 43486 50430 43538
rect 50482 43486 50494 43538
rect 51874 43486 51886 43538
rect 51938 43486 51950 43538
rect 53554 43486 53566 43538
rect 53618 43486 53630 43538
rect 58482 43486 58494 43538
rect 58546 43486 58558 43538
rect 50766 43474 50818 43486
rect 58942 43474 58994 43486
rect 60286 43538 60338 43550
rect 62302 43538 62354 43550
rect 61954 43486 61966 43538
rect 62018 43486 62030 43538
rect 60286 43474 60338 43486
rect 62302 43474 62354 43486
rect 62414 43538 62466 43550
rect 62414 43474 62466 43486
rect 62750 43538 62802 43550
rect 62750 43474 62802 43486
rect 65326 43538 65378 43550
rect 87266 43486 87278 43538
rect 87330 43486 87342 43538
rect 65326 43474 65378 43486
rect 48302 43426 48354 43438
rect 48302 43362 48354 43374
rect 48862 43426 48914 43438
rect 48862 43362 48914 43374
rect 49870 43426 49922 43438
rect 52446 43426 52498 43438
rect 58046 43426 58098 43438
rect 51986 43374 51998 43426
rect 52050 43374 52062 43426
rect 56354 43374 56366 43426
rect 56418 43374 56430 43426
rect 49870 43362 49922 43374
rect 52446 43362 52498 43374
rect 58046 43362 58098 43374
rect 63982 43426 64034 43438
rect 87838 43426 87890 43438
rect 116846 43426 116898 43438
rect 82338 43374 82350 43426
rect 82402 43374 82414 43426
rect 114930 43374 114942 43426
rect 114994 43374 115006 43426
rect 63982 43362 64034 43374
rect 87838 43362 87890 43374
rect 116846 43362 116898 43374
rect 59950 43314 60002 43326
rect 59950 43250 60002 43262
rect 60062 43314 60114 43326
rect 60062 43250 60114 43262
rect 60510 43314 60562 43326
rect 60510 43250 60562 43262
rect 1344 43146 118608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 118608 43146
rect 1344 43060 118608 43094
rect 50430 42866 50482 42878
rect 48738 42814 48750 42866
rect 48802 42814 48814 42866
rect 50430 42802 50482 42814
rect 50878 42866 50930 42878
rect 50878 42802 50930 42814
rect 52222 42866 52274 42878
rect 52222 42802 52274 42814
rect 54910 42866 54962 42878
rect 54910 42802 54962 42814
rect 55358 42866 55410 42878
rect 55358 42802 55410 42814
rect 55918 42866 55970 42878
rect 55918 42802 55970 42814
rect 56366 42866 56418 42878
rect 56366 42802 56418 42814
rect 56702 42866 56754 42878
rect 56702 42802 56754 42814
rect 57262 42866 57314 42878
rect 57262 42802 57314 42814
rect 58830 42866 58882 42878
rect 58830 42802 58882 42814
rect 60622 42866 60674 42878
rect 62190 42866 62242 42878
rect 61730 42814 61742 42866
rect 61794 42814 61806 42866
rect 60622 42802 60674 42814
rect 62190 42802 62242 42814
rect 62750 42866 62802 42878
rect 62750 42802 62802 42814
rect 63198 42866 63250 42878
rect 63198 42802 63250 42814
rect 64430 42866 64482 42878
rect 64430 42802 64482 42814
rect 48190 42754 48242 42766
rect 49870 42754 49922 42766
rect 49522 42702 49534 42754
rect 49586 42702 49598 42754
rect 48190 42690 48242 42702
rect 49870 42690 49922 42702
rect 50206 42754 50258 42766
rect 50206 42690 50258 42702
rect 51550 42754 51602 42766
rect 52558 42754 52610 42766
rect 51762 42702 51774 42754
rect 51826 42702 51838 42754
rect 52098 42702 52110 42754
rect 52162 42702 52174 42754
rect 51550 42690 51602 42702
rect 52558 42690 52610 42702
rect 57934 42754 57986 42766
rect 57934 42690 57986 42702
rect 58270 42754 58322 42766
rect 58270 42690 58322 42702
rect 59166 42754 59218 42766
rect 59166 42690 59218 42702
rect 59614 42754 59666 42766
rect 59614 42690 59666 42702
rect 59950 42754 60002 42766
rect 59950 42690 60002 42702
rect 48974 42642 49026 42654
rect 48974 42578 49026 42590
rect 49758 42642 49810 42654
rect 49758 42578 49810 42590
rect 53454 42642 53506 42654
rect 53454 42578 53506 42590
rect 53678 42642 53730 42654
rect 53678 42578 53730 42590
rect 54238 42642 54290 42654
rect 54238 42578 54290 42590
rect 57710 42642 57762 42654
rect 57710 42578 57762 42590
rect 59502 42642 59554 42654
rect 59502 42578 59554 42590
rect 61406 42642 61458 42654
rect 61406 42578 61458 42590
rect 61630 42642 61682 42654
rect 61630 42578 61682 42590
rect 63534 42642 63586 42654
rect 63534 42578 63586 42590
rect 63982 42642 64034 42654
rect 63982 42578 64034 42590
rect 47742 42530 47794 42542
rect 47742 42466 47794 42478
rect 50542 42530 50594 42542
rect 50542 42466 50594 42478
rect 51438 42530 51490 42542
rect 51438 42466 51490 42478
rect 52670 42530 52722 42542
rect 52670 42466 52722 42478
rect 53566 42530 53618 42542
rect 53566 42466 53618 42478
rect 58046 42530 58098 42542
rect 58046 42466 58098 42478
rect 58158 42530 58210 42542
rect 58158 42466 58210 42478
rect 59390 42530 59442 42542
rect 59390 42466 59442 42478
rect 60062 42530 60114 42542
rect 60062 42466 60114 42478
rect 1344 42362 118608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 118608 42362
rect 1344 42276 118608 42310
rect 56814 42194 56866 42206
rect 63970 42142 63982 42194
rect 64034 42142 64046 42194
rect 56814 42130 56866 42142
rect 58158 42082 58210 42094
rect 61730 42030 61742 42082
rect 61794 42030 61806 42082
rect 58158 42018 58210 42030
rect 55246 41970 55298 41982
rect 54786 41918 54798 41970
rect 54850 41918 54862 41970
rect 55246 41906 55298 41918
rect 55694 41970 55746 41982
rect 114382 41970 114434 41982
rect 57922 41918 57934 41970
rect 57986 41918 57998 41970
rect 59378 41918 59390 41970
rect 59442 41918 59454 41970
rect 60946 41918 60958 41970
rect 61010 41918 61022 41970
rect 114930 41918 114942 41970
rect 114994 41918 115006 41970
rect 55694 41906 55746 41918
rect 114382 41906 114434 41918
rect 48302 41858 48354 41870
rect 48302 41794 48354 41806
rect 48750 41858 48802 41870
rect 57374 41858 57426 41870
rect 60398 41858 60450 41870
rect 52770 41806 52782 41858
rect 52834 41806 52846 41858
rect 59266 41806 59278 41858
rect 59330 41806 59342 41858
rect 115826 41806 115838 41858
rect 115890 41806 115902 41858
rect 48750 41794 48802 41806
rect 57374 41794 57426 41806
rect 60398 41794 60450 41806
rect 58270 41746 58322 41758
rect 59490 41694 59502 41746
rect 59554 41694 59566 41746
rect 60050 41694 60062 41746
rect 60114 41743 60126 41746
rect 60386 41743 60398 41746
rect 60114 41697 60398 41743
rect 60114 41694 60126 41697
rect 60386 41694 60398 41697
rect 60450 41694 60462 41746
rect 58270 41682 58322 41694
rect 1344 41578 118608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 118608 41578
rect 1344 41492 118608 41526
rect 57138 41358 57150 41410
rect 57202 41407 57214 41410
rect 57698 41407 57710 41410
rect 57202 41361 57710 41407
rect 57202 41358 57214 41361
rect 57698 41358 57710 41361
rect 57762 41358 57774 41410
rect 49198 41298 49250 41310
rect 57150 41298 57202 41310
rect 3266 41246 3278 41298
rect 3330 41246 3342 41298
rect 52658 41246 52670 41298
rect 52722 41246 52734 41298
rect 54226 41246 54238 41298
rect 54290 41246 54302 41298
rect 56354 41246 56366 41298
rect 56418 41246 56430 41298
rect 49198 41234 49250 41246
rect 57150 41234 57202 41246
rect 58718 41298 58770 41310
rect 58718 41234 58770 41246
rect 59502 41298 59554 41310
rect 59502 41234 59554 41246
rect 61406 41298 61458 41310
rect 61406 41234 61458 41246
rect 61518 41298 61570 41310
rect 115490 41246 115502 41298
rect 115554 41246 115566 41298
rect 61518 41234 61570 41246
rect 59054 41186 59106 41198
rect 47506 41134 47518 41186
rect 47570 41134 47582 41186
rect 49858 41134 49870 41186
rect 49922 41134 49934 41186
rect 53442 41134 53454 41186
rect 53506 41134 53518 41186
rect 116162 41134 116174 41186
rect 116226 41134 116238 41186
rect 59054 41122 59106 41134
rect 1922 41022 1934 41074
rect 1986 41022 1998 41074
rect 50530 41022 50542 41074
rect 50594 41022 50606 41074
rect 47742 40962 47794 40974
rect 47742 40898 47794 40910
rect 57598 40962 57650 40974
rect 57598 40898 57650 40910
rect 58158 40962 58210 40974
rect 58158 40898 58210 40910
rect 60174 40962 60226 40974
rect 60174 40898 60226 40910
rect 60622 40962 60674 40974
rect 60622 40898 60674 40910
rect 61630 40962 61682 40974
rect 61630 40898 61682 40910
rect 62190 40962 62242 40974
rect 62190 40898 62242 40910
rect 62750 40962 62802 40974
rect 62750 40898 62802 40910
rect 116958 40962 117010 40974
rect 116958 40898 117010 40910
rect 1344 40794 118608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 118608 40794
rect 1344 40708 118608 40742
rect 49422 40626 49474 40638
rect 49422 40562 49474 40574
rect 50878 40626 50930 40638
rect 50878 40562 50930 40574
rect 51550 40626 51602 40638
rect 51550 40562 51602 40574
rect 52334 40626 52386 40638
rect 52334 40562 52386 40574
rect 53118 40626 53170 40638
rect 53118 40562 53170 40574
rect 54126 40626 54178 40638
rect 54126 40562 54178 40574
rect 54462 40626 54514 40638
rect 54462 40562 54514 40574
rect 61966 40626 62018 40638
rect 61966 40562 62018 40574
rect 117070 40626 117122 40638
rect 117070 40562 117122 40574
rect 1710 40514 1762 40526
rect 53678 40514 53730 40526
rect 47954 40462 47966 40514
rect 48018 40462 48030 40514
rect 1710 40450 1762 40462
rect 53678 40450 53730 40462
rect 61182 40514 61234 40526
rect 116274 40462 116286 40514
rect 116338 40462 116350 40514
rect 61182 40450 61234 40462
rect 52670 40402 52722 40414
rect 62414 40402 62466 40414
rect 48738 40350 48750 40402
rect 48802 40350 48814 40402
rect 61506 40350 61518 40402
rect 61570 40350 61582 40402
rect 117282 40350 117294 40402
rect 117346 40350 117358 40402
rect 52670 40338 52722 40350
rect 62414 40338 62466 40350
rect 50654 40290 50706 40302
rect 61294 40290 61346 40302
rect 45826 40238 45838 40290
rect 45890 40238 45902 40290
rect 50978 40238 50990 40290
rect 51042 40238 51054 40290
rect 115154 40238 115166 40290
rect 115218 40238 115230 40290
rect 50654 40226 50706 40238
rect 61294 40226 61346 40238
rect 1344 40010 118608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 118608 40010
rect 1344 39924 118608 39958
rect 48078 39842 48130 39854
rect 48078 39778 48130 39790
rect 3614 39730 3666 39742
rect 3614 39666 3666 39678
rect 47406 39730 47458 39742
rect 47406 39666 47458 39678
rect 48414 39730 48466 39742
rect 48414 39666 48466 39678
rect 49870 39730 49922 39742
rect 49870 39666 49922 39678
rect 51326 39730 51378 39742
rect 51326 39666 51378 39678
rect 53342 39730 53394 39742
rect 53342 39666 53394 39678
rect 117070 39730 117122 39742
rect 117070 39666 117122 39678
rect 3042 39566 3054 39618
rect 3106 39566 3118 39618
rect 49186 39566 49198 39618
rect 49250 39566 49262 39618
rect 50206 39506 50258 39518
rect 1922 39454 1934 39506
rect 1986 39454 1998 39506
rect 48962 39454 48974 39506
rect 49026 39454 49038 39506
rect 50206 39442 50258 39454
rect 1344 39226 118608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 118608 39226
rect 1344 39140 118608 39174
rect 61070 39058 61122 39070
rect 61070 38994 61122 39006
rect 63422 39058 63474 39070
rect 63422 38994 63474 39006
rect 53790 38946 53842 38958
rect 63870 38946 63922 38958
rect 62850 38894 62862 38946
rect 62914 38894 62926 38946
rect 53790 38882 53842 38894
rect 63870 38882 63922 38894
rect 118078 38946 118130 38958
rect 118078 38882 118130 38894
rect 62078 38834 62130 38846
rect 53554 38782 53566 38834
rect 53618 38782 53630 38834
rect 62626 38782 62638 38834
rect 62690 38782 62702 38834
rect 62078 38770 62130 38782
rect 61742 38610 61794 38622
rect 61742 38546 61794 38558
rect 1344 38442 118608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 118608 38442
rect 1344 38356 118608 38390
rect 52782 38162 52834 38174
rect 54226 38110 54238 38162
rect 54290 38110 54302 38162
rect 56354 38110 56366 38162
rect 56418 38110 56430 38162
rect 64306 38110 64318 38162
rect 64370 38110 64382 38162
rect 52782 38098 52834 38110
rect 3042 37998 3054 38050
rect 3106 37998 3118 38050
rect 53442 37998 53454 38050
rect 53506 37998 53518 38050
rect 61394 37998 61406 38050
rect 61458 37998 61470 38050
rect 1922 37886 1934 37938
rect 1986 37886 1998 37938
rect 62178 37886 62190 37938
rect 62242 37886 62254 37938
rect 3502 37826 3554 37838
rect 3502 37762 3554 37774
rect 60622 37826 60674 37838
rect 60622 37762 60674 37774
rect 1344 37658 118608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 118608 37658
rect 1344 37572 118608 37606
rect 54238 37490 54290 37502
rect 54238 37426 54290 37438
rect 56030 37490 56082 37502
rect 56030 37426 56082 37438
rect 61854 37490 61906 37502
rect 61854 37426 61906 37438
rect 1922 37326 1934 37378
rect 1986 37326 1998 37378
rect 54898 37326 54910 37378
rect 54962 37326 54974 37378
rect 55122 37326 55134 37378
rect 55186 37326 55198 37378
rect 54574 37266 54626 37278
rect 61618 37214 61630 37266
rect 61682 37214 61694 37266
rect 54574 37202 54626 37214
rect 53566 37154 53618 37166
rect 3266 37102 3278 37154
rect 3330 37102 3342 37154
rect 53566 37090 53618 37102
rect 56366 37154 56418 37166
rect 56366 37090 56418 37102
rect 1344 36874 118608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 118608 36874
rect 1344 36788 118608 36822
rect 3266 36542 3278 36594
rect 3330 36542 3342 36594
rect 114818 36542 114830 36594
rect 114882 36542 114894 36594
rect 2146 36318 2158 36370
rect 2210 36318 2222 36370
rect 116162 36318 116174 36370
rect 116226 36318 116238 36370
rect 117070 36258 117122 36270
rect 117070 36194 117122 36206
rect 1344 36090 118608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 118608 36090
rect 1344 36004 118608 36038
rect 1822 35922 1874 35934
rect 1822 35858 1874 35870
rect 2158 35810 2210 35822
rect 2158 35746 2210 35758
rect 114494 35698 114546 35710
rect 114930 35646 114942 35698
rect 114994 35646 115006 35698
rect 114494 35634 114546 35646
rect 115826 35534 115838 35586
rect 115890 35534 115902 35586
rect 1344 35306 118608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 118608 35306
rect 1344 35220 118608 35254
rect 3266 34974 3278 35026
rect 3330 34974 3342 35026
rect 45826 34862 45838 34914
rect 45890 34862 45902 34914
rect 116162 34862 116174 34914
rect 116226 34862 116238 34914
rect 58270 34802 58322 34814
rect 1922 34750 1934 34802
rect 1986 34750 1998 34802
rect 58270 34738 58322 34750
rect 46062 34690 46114 34702
rect 46062 34626 46114 34638
rect 57710 34690 57762 34702
rect 57710 34626 57762 34638
rect 58606 34690 58658 34702
rect 58606 34626 58658 34638
rect 115950 34690 116002 34702
rect 115950 34626 116002 34638
rect 1344 34522 118608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 118608 34522
rect 1344 34436 118608 34470
rect 47170 34190 47182 34242
rect 47234 34190 47246 34242
rect 115938 34190 115950 34242
rect 116002 34190 116014 34242
rect 3042 34078 3054 34130
rect 3106 34078 3118 34130
rect 47954 34078 47966 34130
rect 48018 34078 48030 34130
rect 115154 34078 115166 34130
rect 115218 34078 115230 34130
rect 3614 34018 3666 34030
rect 48414 34018 48466 34030
rect 1922 33966 1934 34018
rect 1986 33966 1998 34018
rect 45042 33966 45054 34018
rect 45106 33966 45118 34018
rect 3614 33954 3666 33966
rect 48414 33954 48466 33966
rect 114606 34018 114658 34030
rect 118066 33966 118078 34018
rect 118130 33966 118142 34018
rect 114606 33954 114658 33966
rect 1344 33738 118608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 118608 33738
rect 1344 33652 118608 33686
rect 46062 33570 46114 33582
rect 46062 33506 46114 33518
rect 1822 33458 1874 33470
rect 1822 33394 1874 33406
rect 45390 33458 45442 33470
rect 45390 33394 45442 33406
rect 46398 33458 46450 33470
rect 46398 33394 46450 33406
rect 47742 33458 47794 33470
rect 115490 33406 115502 33458
rect 115554 33406 115566 33458
rect 47742 33394 47794 33406
rect 48190 33346 48242 33358
rect 116050 33294 116062 33346
rect 116114 33294 116126 33346
rect 48190 33282 48242 33294
rect 46610 33182 46622 33234
rect 46674 33182 46686 33234
rect 46946 33182 46958 33234
rect 47010 33182 47022 33234
rect 1344 32954 118608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 118608 32954
rect 1344 32868 118608 32902
rect 116062 32786 116114 32798
rect 116062 32722 116114 32734
rect 114942 32674 114994 32686
rect 1922 32622 1934 32674
rect 1986 32622 1998 32674
rect 116610 32622 116622 32674
rect 116674 32622 116686 32674
rect 117170 32622 117182 32674
rect 117234 32622 117246 32674
rect 114942 32610 114994 32622
rect 115390 32450 115442 32462
rect 3266 32398 3278 32450
rect 3330 32398 3342 32450
rect 115390 32386 115442 32398
rect 116398 32338 116450 32350
rect 116398 32274 116450 32286
rect 1344 32170 118608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 118608 32170
rect 1344 32084 118608 32118
rect 1822 31890 1874 31902
rect 1822 31826 1874 31838
rect 1344 31386 118608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 118608 31386
rect 1344 31300 118608 31334
rect 116162 30942 116174 30994
rect 116226 30942 116238 30994
rect 115490 30830 115502 30882
rect 115554 30830 115566 30882
rect 1344 30602 118608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 118608 30602
rect 1344 30516 118608 30550
rect 116162 30382 116174 30434
rect 116226 30431 116238 30434
rect 116498 30431 116510 30434
rect 116226 30385 116510 30431
rect 116226 30382 116238 30385
rect 116498 30382 116510 30385
rect 116562 30382 116574 30434
rect 3266 30270 3278 30322
rect 3330 30270 3342 30322
rect 114382 30210 114434 30222
rect 69346 30158 69358 30210
rect 69410 30158 69422 30210
rect 114382 30146 114434 30158
rect 114942 30210 114994 30222
rect 114942 30146 114994 30158
rect 115502 30210 115554 30222
rect 115502 30146 115554 30158
rect 117070 30098 117122 30110
rect 1922 30046 1934 30098
rect 1986 30046 1998 30098
rect 72258 30046 72270 30098
rect 72322 30046 72334 30098
rect 117070 30034 117122 30046
rect 117406 30098 117458 30110
rect 117406 30034 117458 30046
rect 75070 29986 75122 29998
rect 75070 29922 75122 29934
rect 116286 29986 116338 29998
rect 116286 29922 116338 29934
rect 1344 29818 118608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 118608 29818
rect 1344 29732 118608 29766
rect 1822 29650 1874 29662
rect 1822 29586 1874 29598
rect 49422 29650 49474 29662
rect 49422 29586 49474 29598
rect 47730 29374 47742 29426
rect 47794 29374 47806 29426
rect 48526 29202 48578 29214
rect 48526 29138 48578 29150
rect 1344 29034 118608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 118608 29034
rect 1344 28948 118608 28982
rect 45502 28530 45554 28542
rect 45502 28466 45554 28478
rect 45838 28418 45890 28430
rect 45838 28354 45890 28366
rect 1344 28250 118608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 118608 28250
rect 1344 28164 118608 28198
rect 48190 28082 48242 28094
rect 48190 28018 48242 28030
rect 46946 27918 46958 27970
rect 47010 27918 47022 27970
rect 47730 27806 47742 27858
rect 47794 27806 47806 27858
rect 44818 27694 44830 27746
rect 44882 27694 44894 27746
rect 1344 27466 118608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 118608 27466
rect 1344 27380 118608 27414
rect 45726 27298 45778 27310
rect 45726 27234 45778 27246
rect 46062 27298 46114 27310
rect 46062 27234 46114 27246
rect 47406 27186 47458 27198
rect 3266 27134 3278 27186
rect 3330 27134 3342 27186
rect 47406 27122 47458 27134
rect 47854 27186 47906 27198
rect 115490 27134 115502 27186
rect 115554 27134 115566 27186
rect 47854 27122 47906 27134
rect 46834 27022 46846 27074
rect 46898 27022 46910 27074
rect 116162 27022 116174 27074
rect 116226 27022 116238 27074
rect 44718 26962 44770 26974
rect 117070 26962 117122 26974
rect 1922 26910 1934 26962
rect 1986 26910 1998 26962
rect 46610 26910 46622 26962
rect 46674 26910 46686 26962
rect 44718 26898 44770 26910
rect 117070 26898 117122 26910
rect 117406 26962 117458 26974
rect 117406 26898 117458 26910
rect 1344 26682 118608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 118608 26682
rect 1344 26596 118608 26630
rect 63198 26514 63250 26526
rect 63198 26450 63250 26462
rect 116734 26514 116786 26526
rect 116734 26450 116786 26462
rect 1710 26402 1762 26414
rect 58818 26350 58830 26402
rect 58882 26350 58894 26402
rect 1710 26338 1762 26350
rect 114382 26290 114434 26302
rect 62738 26238 62750 26290
rect 62802 26238 62814 26290
rect 114930 26238 114942 26290
rect 114994 26238 115006 26290
rect 114382 26226 114434 26238
rect 2158 26178 2210 26190
rect 115826 26126 115838 26178
rect 115890 26126 115902 26178
rect 2158 26114 2210 26126
rect 1344 25898 118608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 118608 25898
rect 1344 25812 118608 25846
rect 3266 25566 3278 25618
rect 3330 25566 3342 25618
rect 45602 25454 45614 25506
rect 45666 25454 45678 25506
rect 1922 25342 1934 25394
rect 1986 25342 1998 25394
rect 45838 25282 45890 25294
rect 45838 25218 45890 25230
rect 1344 25114 118608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 118608 25114
rect 1344 25028 118608 25062
rect 48078 24946 48130 24958
rect 48078 24882 48130 24894
rect 46834 24782 46846 24834
rect 46898 24782 46910 24834
rect 3042 24670 3054 24722
rect 3106 24670 3118 24722
rect 47618 24670 47630 24722
rect 47682 24670 47694 24722
rect 3502 24610 3554 24622
rect 1922 24558 1934 24610
rect 1986 24558 1998 24610
rect 44706 24558 44718 24610
rect 44770 24558 44782 24610
rect 3502 24546 3554 24558
rect 1344 24330 118608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 118608 24330
rect 1344 24244 118608 24278
rect 45726 24162 45778 24174
rect 77858 24110 77870 24162
rect 77922 24159 77934 24162
rect 78418 24159 78430 24162
rect 77922 24113 78430 24159
rect 77922 24110 77934 24113
rect 78418 24110 78430 24113
rect 78482 24110 78494 24162
rect 45726 24098 45778 24110
rect 77870 24050 77922 24062
rect 77870 23986 77922 23998
rect 46062 23938 46114 23950
rect 46834 23886 46846 23938
rect 46898 23886 46910 23938
rect 46062 23874 46114 23886
rect 44718 23826 44770 23838
rect 47406 23826 47458 23838
rect 46610 23774 46622 23826
rect 46674 23774 46686 23826
rect 44718 23762 44770 23774
rect 47406 23762 47458 23774
rect 47854 23714 47906 23726
rect 47854 23650 47906 23662
rect 78318 23714 78370 23726
rect 78318 23650 78370 23662
rect 1344 23546 118608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 118608 23546
rect 1344 23460 118608 23494
rect 116622 23378 116674 23390
rect 116622 23314 116674 23326
rect 45838 23266 45890 23278
rect 45838 23202 45890 23214
rect 77870 23266 77922 23278
rect 117070 23266 117122 23278
rect 79090 23214 79102 23266
rect 79154 23214 79166 23266
rect 79650 23214 79662 23266
rect 79714 23214 79726 23266
rect 77870 23202 77922 23214
rect 117070 23202 117122 23214
rect 78542 23154 78594 23166
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 45602 23102 45614 23154
rect 45666 23102 45678 23154
rect 77634 23102 77646 23154
rect 77698 23102 77710 23154
rect 78542 23090 78594 23102
rect 78878 23154 78930 23166
rect 117282 23102 117294 23154
rect 117346 23102 117358 23154
rect 78878 23090 78930 23102
rect 3502 23042 3554 23054
rect 1922 22990 1934 23042
rect 1986 22990 1998 23042
rect 3502 22978 3554 22990
rect 80222 23042 80274 23054
rect 80222 22978 80274 22990
rect 1344 22762 118608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 118608 22762
rect 1344 22676 118608 22710
rect 48190 22482 48242 22494
rect 48190 22418 48242 22430
rect 76526 22482 76578 22494
rect 78306 22430 78318 22482
rect 78370 22430 78382 22482
rect 80434 22430 80446 22482
rect 80498 22430 80510 22482
rect 115490 22430 115502 22482
rect 115554 22430 115566 22482
rect 76526 22418 76578 22430
rect 46398 22370 46450 22382
rect 47170 22318 47182 22370
rect 47234 22318 47246 22370
rect 77522 22318 77534 22370
rect 77586 22318 77598 22370
rect 116162 22318 116174 22370
rect 116226 22318 116238 22370
rect 46398 22306 46450 22318
rect 47742 22258 47794 22270
rect 1922 22206 1934 22258
rect 1986 22206 1998 22258
rect 46946 22206 46958 22258
rect 47010 22206 47022 22258
rect 47742 22194 47794 22206
rect 91758 22258 91810 22270
rect 91758 22194 91810 22206
rect 4398 22146 4450 22158
rect 4398 22082 4450 22094
rect 45502 22146 45554 22158
rect 45502 22082 45554 22094
rect 46062 22146 46114 22158
rect 46062 22082 46114 22094
rect 92094 22146 92146 22158
rect 92094 22082 92146 22094
rect 1344 21978 118608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 118608 21978
rect 1344 21892 118608 21926
rect 48414 21810 48466 21822
rect 48414 21746 48466 21758
rect 44494 21698 44546 21710
rect 47170 21646 47182 21698
rect 47234 21646 47246 21698
rect 91970 21646 91982 21698
rect 92034 21646 92046 21698
rect 44494 21634 44546 21646
rect 3042 21534 3054 21586
rect 3106 21534 3118 21586
rect 44258 21534 44270 21586
rect 44322 21534 44334 21586
rect 47954 21534 47966 21586
rect 48018 21534 48030 21586
rect 91298 21534 91310 21586
rect 91362 21534 91374 21586
rect 3614 21474 3666 21486
rect 90638 21474 90690 21486
rect 1922 21422 1934 21474
rect 1986 21422 1998 21474
rect 45042 21422 45054 21474
rect 45106 21422 45118 21474
rect 94098 21422 94110 21474
rect 94162 21422 94174 21474
rect 3614 21410 3666 21422
rect 90638 21410 90690 21422
rect 1344 21194 118608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 118608 21194
rect 1344 21108 118608 21142
rect 91198 21026 91250 21038
rect 91198 20962 91250 20974
rect 1822 20914 1874 20926
rect 1822 20850 1874 20862
rect 40238 20914 40290 20926
rect 48974 20914 49026 20926
rect 45490 20862 45502 20914
rect 45554 20862 45566 20914
rect 47618 20862 47630 20914
rect 47682 20862 47694 20914
rect 40238 20850 40290 20862
rect 48974 20850 49026 20862
rect 93102 20914 93154 20926
rect 93102 20850 93154 20862
rect 39790 20802 39842 20814
rect 91534 20802 91586 20814
rect 48290 20750 48302 20802
rect 48354 20750 48366 20802
rect 92194 20750 92206 20802
rect 92258 20750 92270 20802
rect 39790 20738 39842 20750
rect 91534 20738 91586 20750
rect 39454 20690 39506 20702
rect 92306 20638 92318 20690
rect 92370 20638 92382 20690
rect 39454 20626 39506 20638
rect 90078 20578 90130 20590
rect 90078 20514 90130 20526
rect 90526 20578 90578 20590
rect 90526 20514 90578 20526
rect 1344 20410 118608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 118608 20410
rect 1344 20324 118608 20358
rect 45502 20130 45554 20142
rect 45502 20066 45554 20078
rect 46062 20130 46114 20142
rect 46946 20078 46958 20130
rect 47010 20078 47022 20130
rect 46062 20066 46114 20078
rect 48302 20018 48354 20030
rect 47170 19966 47182 20018
rect 47234 19966 47246 20018
rect 48302 19954 48354 19966
rect 47742 19906 47794 19918
rect 47742 19842 47794 19854
rect 46398 19794 46450 19806
rect 46398 19730 46450 19742
rect 1344 19626 118608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 118608 19626
rect 1344 19540 118608 19574
rect 115490 19294 115502 19346
rect 115554 19294 115566 19346
rect 117406 19234 117458 19246
rect 116162 19182 116174 19234
rect 116226 19182 116238 19234
rect 117406 19170 117458 19182
rect 117070 19122 117122 19134
rect 117070 19058 117122 19070
rect 1344 18842 118608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 118608 18842
rect 1344 18756 118608 18790
rect 116734 18674 116786 18686
rect 116734 18610 116786 18622
rect 1822 18562 1874 18574
rect 1822 18498 1874 18510
rect 1344 18058 118608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 118608 18058
rect 1344 17972 118608 18006
rect 1822 17442 1874 17454
rect 1822 17378 1874 17390
rect 1344 17274 118608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 118608 17274
rect 1344 17188 118608 17222
rect 118078 16994 118130 17006
rect 118078 16930 118130 16942
rect 3502 16882 3554 16894
rect 3042 16830 3054 16882
rect 3106 16830 3118 16882
rect 3502 16818 3554 16830
rect 1922 16718 1934 16770
rect 1986 16718 1998 16770
rect 1344 16490 118608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 118608 16490
rect 1344 16404 118608 16438
rect 1344 15706 118608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 118608 15706
rect 1344 15620 118608 15654
rect 54462 15426 54514 15438
rect 54462 15362 54514 15374
rect 114494 15426 114546 15438
rect 114494 15362 114546 15374
rect 54126 15314 54178 15326
rect 114930 15262 114942 15314
rect 114994 15262 115006 15314
rect 54126 15250 54178 15262
rect 53678 15202 53730 15214
rect 115826 15150 115838 15202
rect 115890 15150 115902 15202
rect 53678 15138 53730 15150
rect 1344 14922 118608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 118608 14922
rect 1344 14836 118608 14870
rect 115826 14590 115838 14642
rect 115890 14590 115902 14642
rect 114494 14530 114546 14542
rect 114930 14478 114942 14530
rect 114994 14478 115006 14530
rect 114494 14466 114546 14478
rect 1344 14138 118608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 118608 14138
rect 1344 14052 118608 14086
rect 1344 13354 118608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 118608 13354
rect 1344 13268 118608 13302
rect 1344 12570 118608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 118608 12570
rect 1344 12484 118608 12518
rect 116274 12238 116286 12290
rect 116338 12238 116350 12290
rect 2818 12126 2830 12178
rect 2882 12126 2894 12178
rect 116846 12066 116898 12078
rect 1922 12014 1934 12066
rect 1986 12014 1998 12066
rect 114930 12014 114942 12066
rect 114994 12014 115006 12066
rect 116846 12002 116898 12014
rect 1344 11786 118608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 118608 11786
rect 1344 11700 118608 11734
rect 3278 11506 3330 11518
rect 3278 11442 3330 11454
rect 2594 11342 2606 11394
rect 2658 11342 2670 11394
rect 2830 11282 2882 11294
rect 2830 11218 2882 11230
rect 1344 11002 118608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 118608 11002
rect 1344 10916 118608 10950
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 3502 10498 3554 10510
rect 1922 10446 1934 10498
rect 1986 10446 1998 10498
rect 3502 10434 3554 10446
rect 1344 10218 118608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 118608 10218
rect 1344 10132 118608 10166
rect 115490 9886 115502 9938
rect 115554 9886 115566 9938
rect 116162 9774 116174 9826
rect 116226 9774 116238 9826
rect 117282 9774 117294 9826
rect 117346 9774 117358 9826
rect 117070 9714 117122 9726
rect 117070 9650 117122 9662
rect 1344 9434 118608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 118608 9434
rect 1344 9348 118608 9382
rect 116734 9266 116786 9278
rect 116734 9202 116786 9214
rect 1344 8650 118608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 118608 8650
rect 1344 8564 118608 8598
rect 63870 8370 63922 8382
rect 115826 8318 115838 8370
rect 115890 8318 115902 8370
rect 63870 8306 63922 8318
rect 64430 8258 64482 8270
rect 64430 8194 64482 8206
rect 114494 8258 114546 8270
rect 114930 8206 114942 8258
rect 114994 8206 115006 8258
rect 114494 8194 114546 8206
rect 64766 8034 64818 8046
rect 64766 7970 64818 7982
rect 1344 7866 118608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 118608 7866
rect 1344 7780 118608 7814
rect 1822 7586 1874 7598
rect 1822 7522 1874 7534
rect 116162 7422 116174 7474
rect 116226 7422 116238 7474
rect 2382 7362 2434 7374
rect 116734 7362 116786 7374
rect 115490 7310 115502 7362
rect 115554 7310 115566 7362
rect 2382 7298 2434 7310
rect 116734 7298 116786 7310
rect 1344 7082 118608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 118608 7082
rect 1344 6996 118608 7030
rect 114818 6750 114830 6802
rect 114882 6750 114894 6802
rect 3042 6638 3054 6690
rect 3106 6638 3118 6690
rect 117070 6578 117122 6590
rect 1922 6526 1934 6578
rect 1986 6526 1998 6578
rect 116162 6526 116174 6578
rect 116226 6526 116238 6578
rect 117070 6514 117122 6526
rect 117406 6578 117458 6590
rect 117406 6514 117458 6526
rect 3614 6466 3666 6478
rect 3614 6402 3666 6414
rect 1344 6298 118608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 118608 6298
rect 1344 6212 118608 6246
rect 112366 6130 112418 6142
rect 112366 6066 112418 6078
rect 116274 5966 116286 6018
rect 116338 5966 116350 6018
rect 3502 5906 3554 5918
rect 3042 5854 3054 5906
rect 3106 5854 3118 5906
rect 113138 5854 113150 5906
rect 113202 5854 113214 5906
rect 3502 5842 3554 5854
rect 5182 5794 5234 5806
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 5182 5730 5234 5742
rect 42030 5794 42082 5806
rect 42030 5730 42082 5742
rect 48078 5794 48130 5806
rect 116846 5794 116898 5806
rect 113810 5742 113822 5794
rect 113874 5742 113886 5794
rect 114930 5742 114942 5794
rect 114994 5742 115006 5794
rect 48078 5730 48130 5742
rect 116846 5730 116898 5742
rect 117294 5794 117346 5806
rect 117294 5730 117346 5742
rect 1344 5514 118608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 118608 5514
rect 1344 5428 118608 5462
rect 5630 5234 5682 5246
rect 5630 5170 5682 5182
rect 6078 5234 6130 5246
rect 6078 5170 6130 5182
rect 43262 5234 43314 5246
rect 43262 5170 43314 5182
rect 46174 5234 46226 5246
rect 49198 5234 49250 5246
rect 47282 5182 47294 5234
rect 47346 5182 47358 5234
rect 46174 5170 46226 5182
rect 49198 5170 49250 5182
rect 50318 5234 50370 5246
rect 112802 5182 112814 5234
rect 112866 5182 112878 5234
rect 114818 5182 114830 5234
rect 114882 5182 114894 5234
rect 50318 5170 50370 5182
rect 25230 5122 25282 5134
rect 26910 5122 26962 5134
rect 59838 5122 59890 5134
rect 2818 5070 2830 5122
rect 2882 5070 2894 5122
rect 4834 5070 4846 5122
rect 4898 5070 4910 5122
rect 26338 5070 26350 5122
rect 26402 5070 26414 5122
rect 41570 5070 41582 5122
rect 41634 5070 41646 5122
rect 46610 5070 46622 5122
rect 46674 5070 46686 5122
rect 25230 5058 25282 5070
rect 26910 5058 26962 5070
rect 59838 5058 59890 5070
rect 63982 5122 64034 5134
rect 63982 5058 64034 5070
rect 42366 5010 42418 5022
rect 1922 4958 1934 5010
rect 1986 4958 1998 5010
rect 3714 4958 3726 5010
rect 3778 4958 3790 5010
rect 40674 4958 40686 5010
rect 40738 4958 40750 5010
rect 42366 4946 42418 4958
rect 48414 5010 48466 5022
rect 48414 4946 48466 4958
rect 54798 5010 54850 5022
rect 54798 4946 54850 4958
rect 55246 5010 55298 5022
rect 55246 4946 55298 4958
rect 99150 5010 99202 5022
rect 99150 4946 99202 4958
rect 111358 5010 111410 5022
rect 111358 4946 111410 4958
rect 111918 5010 111970 5022
rect 114146 4958 114158 5010
rect 114210 4958 114222 5010
rect 116162 4958 116174 5010
rect 116226 4958 116238 5010
rect 111918 4946 111970 4958
rect 42702 4898 42754 4910
rect 42702 4834 42754 4846
rect 43710 4898 43762 4910
rect 43710 4834 43762 4846
rect 48750 4898 48802 4910
rect 48750 4834 48802 4846
rect 54462 4898 54514 4910
rect 54462 4834 54514 4846
rect 99486 4898 99538 4910
rect 99486 4834 99538 4846
rect 99934 4898 99986 4910
rect 99934 4834 99986 4846
rect 101390 4898 101442 4910
rect 101390 4834 101442 4846
rect 112254 4898 112306 4910
rect 112254 4834 112306 4846
rect 117070 4898 117122 4910
rect 117070 4834 117122 4846
rect 1344 4730 118608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 118608 4730
rect 1344 4644 118608 4678
rect 6526 4562 6578 4574
rect 6526 4498 6578 4510
rect 9662 4562 9714 4574
rect 9662 4498 9714 4510
rect 10558 4562 10610 4574
rect 10558 4498 10610 4510
rect 11902 4562 11954 4574
rect 11902 4498 11954 4510
rect 15374 4562 15426 4574
rect 15374 4498 15426 4510
rect 28142 4562 28194 4574
rect 28142 4498 28194 4510
rect 32846 4562 32898 4574
rect 32846 4498 32898 4510
rect 46846 4562 46898 4574
rect 46846 4498 46898 4510
rect 49422 4562 49474 4574
rect 49422 4498 49474 4510
rect 57374 4562 57426 4574
rect 57374 4498 57426 4510
rect 62974 4562 63026 4574
rect 62974 4498 63026 4510
rect 65326 4562 65378 4574
rect 65326 4498 65378 4510
rect 68686 4562 68738 4574
rect 68686 4498 68738 4510
rect 76526 4562 76578 4574
rect 76526 4498 76578 4510
rect 78318 4562 78370 4574
rect 78318 4498 78370 4510
rect 80558 4562 80610 4574
rect 80558 4498 80610 4510
rect 81678 4562 81730 4574
rect 81678 4498 81730 4510
rect 104302 4562 104354 4574
rect 104302 4498 104354 4510
rect 5630 4450 5682 4462
rect 1922 4398 1934 4450
rect 1986 4398 1998 4450
rect 5630 4386 5682 4398
rect 5966 4450 6018 4462
rect 5966 4386 6018 4398
rect 11454 4450 11506 4462
rect 45950 4450 46002 4462
rect 18498 4398 18510 4450
rect 18562 4398 18574 4450
rect 44034 4398 44046 4450
rect 44098 4398 44110 4450
rect 11454 4386 11506 4398
rect 45950 4386 46002 4398
rect 46286 4450 46338 4462
rect 46286 4386 46338 4398
rect 49982 4450 50034 4462
rect 49982 4386 50034 4398
rect 50654 4450 50706 4462
rect 50654 4386 50706 4398
rect 50990 4450 51042 4462
rect 67790 4450 67842 4462
rect 53442 4398 53454 4450
rect 53506 4398 53518 4450
rect 61058 4398 61070 4450
rect 61122 4398 61134 4450
rect 50990 4386 51042 4398
rect 67790 4386 67842 4398
rect 68126 4450 68178 4462
rect 76974 4450 77026 4462
rect 71810 4398 71822 4450
rect 71874 4398 71886 4450
rect 68126 4386 68178 4398
rect 76974 4386 77026 4398
rect 77310 4450 77362 4462
rect 101166 4450 101218 4462
rect 87938 4398 87950 4450
rect 88002 4398 88014 4450
rect 93986 4398 93998 4450
rect 94050 4398 94062 4450
rect 99362 4398 99374 4450
rect 99426 4398 99438 4450
rect 77310 4386 77362 4398
rect 101166 4386 101218 4398
rect 103518 4450 103570 4462
rect 103518 4386 103570 4398
rect 103854 4450 103906 4462
rect 117070 4450 117122 4462
rect 116274 4398 116286 4450
rect 116338 4398 116350 4450
rect 103854 4386 103906 4398
rect 117070 4386 117122 4398
rect 117406 4450 117458 4462
rect 117406 4386 117458 4398
rect 4946 4286 4958 4338
rect 5010 4286 5022 4338
rect 8194 4286 8206 4338
rect 8258 4286 8270 4338
rect 11218 4286 11230 4338
rect 11282 4286 11294 4338
rect 14914 4286 14926 4338
rect 14978 4286 14990 4338
rect 27682 4286 27694 4338
rect 27746 4286 27758 4338
rect 32162 4286 32174 4338
rect 32226 4286 32238 4338
rect 43138 4286 43150 4338
rect 43202 4286 43214 4338
rect 48514 4286 48526 4338
rect 48578 4286 48590 4338
rect 51538 4286 51550 4338
rect 51602 4286 51614 4338
rect 56578 4286 56590 4338
rect 56642 4286 56654 4338
rect 59490 4286 59502 4338
rect 59554 4286 59566 4338
rect 63410 4286 63422 4338
rect 63474 4286 63486 4338
rect 73378 4286 73390 4338
rect 73442 4286 73454 4338
rect 78866 4286 78878 4338
rect 78930 4286 78942 4338
rect 83458 4286 83470 4338
rect 83522 4286 83534 4338
rect 94994 4286 95006 4338
rect 95058 4286 95070 4338
rect 100930 4286 100942 4338
rect 100994 4286 101006 4338
rect 101714 4286 101726 4338
rect 101778 4286 101790 4338
rect 112354 4286 112366 4338
rect 112418 4286 112430 4338
rect 113138 4286 113150 4338
rect 113202 4286 113214 4338
rect 8766 4226 8818 4238
rect 17950 4226 18002 4238
rect 21198 4226 21250 4238
rect 3266 4174 3278 4226
rect 3330 4174 3342 4226
rect 3938 4174 3950 4226
rect 4002 4174 4014 4226
rect 7074 4174 7086 4226
rect 7138 4174 7150 4226
rect 13794 4174 13806 4226
rect 13858 4174 13870 4226
rect 19618 4174 19630 4226
rect 19682 4174 19694 4226
rect 8766 4162 8818 4174
rect 17950 4162 18002 4174
rect 21198 4162 21250 4174
rect 21534 4226 21586 4238
rect 36542 4226 36594 4238
rect 26562 4174 26574 4226
rect 26626 4174 26638 4226
rect 31266 4174 31278 4226
rect 31330 4174 31342 4226
rect 21534 4162 21586 4174
rect 36542 4162 36594 4174
rect 37662 4226 37714 4238
rect 70366 4226 70418 4238
rect 75742 4226 75794 4238
rect 86494 4226 86546 4238
rect 92542 4226 92594 4238
rect 97918 4226 97970 4238
rect 100270 4226 100322 4238
rect 117854 4226 117906 4238
rect 42242 4174 42254 4226
rect 42306 4174 42318 4226
rect 45378 4174 45390 4226
rect 45442 4174 45454 4226
rect 47394 4174 47406 4226
rect 47458 4174 47470 4226
rect 52210 4174 52222 4226
rect 52274 4174 52286 4226
rect 54674 4174 54686 4226
rect 54738 4174 54750 4226
rect 55458 4174 55470 4226
rect 55522 4174 55534 4226
rect 58370 4174 58382 4226
rect 58434 4174 58446 4226
rect 60050 4174 60062 4226
rect 60114 4174 60126 4226
rect 64082 4174 64094 4226
rect 64146 4174 64158 4226
rect 70802 4174 70814 4226
rect 70866 4174 70878 4226
rect 74050 4174 74062 4226
rect 74114 4174 74126 4226
rect 79538 4174 79550 4226
rect 79602 4174 79614 4226
rect 82338 4174 82350 4226
rect 82402 4174 82414 4226
rect 86930 4174 86942 4226
rect 86994 4174 87006 4226
rect 92978 4174 92990 4226
rect 93042 4174 93054 4226
rect 95666 4174 95678 4226
rect 95730 4174 95742 4226
rect 98354 4174 98366 4226
rect 98418 4174 98430 4226
rect 102386 4174 102398 4226
rect 102450 4174 102462 4226
rect 111682 4174 111694 4226
rect 111746 4174 111758 4226
rect 113810 4174 113822 4226
rect 113874 4174 113886 4226
rect 114930 4174 114942 4226
rect 114994 4174 115006 4226
rect 37662 4162 37714 4174
rect 70366 4162 70418 4174
rect 75742 4162 75794 4174
rect 86494 4162 86546 4174
rect 92542 4162 92594 4174
rect 97918 4162 97970 4174
rect 100270 4162 100322 4174
rect 117854 4162 117906 4174
rect 1344 3946 118608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 118608 3946
rect 1344 3860 118608 3894
rect 73166 3666 73218 3678
rect 88510 3666 88562 3678
rect 94782 3666 94834 3678
rect 117406 3666 117458 3678
rect 4946 3614 4958 3666
rect 5010 3614 5022 3666
rect 6402 3614 6414 3666
rect 6466 3614 6478 3666
rect 7970 3614 7982 3666
rect 8034 3614 8046 3666
rect 12226 3614 12238 3666
rect 12290 3614 12302 3666
rect 16482 3614 16494 3666
rect 16546 3614 16558 3666
rect 20626 3614 20638 3666
rect 20690 3614 20702 3666
rect 22642 3614 22654 3666
rect 22706 3614 22718 3666
rect 26786 3614 26798 3666
rect 26850 3614 26862 3666
rect 31042 3614 31054 3666
rect 31106 3614 31118 3666
rect 35522 3614 35534 3666
rect 35586 3614 35598 3666
rect 39106 3614 39118 3666
rect 39170 3614 39182 3666
rect 43250 3614 43262 3666
rect 43314 3614 43326 3666
rect 46498 3614 46510 3666
rect 46562 3614 46574 3666
rect 49522 3614 49534 3666
rect 49586 3614 49598 3666
rect 54674 3614 54686 3666
rect 54738 3614 54750 3666
rect 59490 3614 59502 3666
rect 59554 3614 59566 3666
rect 63746 3614 63758 3666
rect 63810 3614 63822 3666
rect 65426 3614 65438 3666
rect 65490 3614 65502 3666
rect 69458 3614 69470 3666
rect 69522 3614 69534 3666
rect 74162 3614 74174 3666
rect 74226 3614 74238 3666
rect 78194 3614 78206 3666
rect 78258 3614 78270 3666
rect 81666 3614 81678 3666
rect 81730 3614 81742 3666
rect 84130 3614 84142 3666
rect 84194 3614 84206 3666
rect 91970 3614 91982 3666
rect 92034 3614 92046 3666
rect 96338 3614 96350 3666
rect 96402 3614 96414 3666
rect 100482 3614 100494 3666
rect 100546 3614 100558 3666
rect 104402 3614 104414 3666
rect 104466 3614 104478 3666
rect 111570 3614 111582 3666
rect 111634 3614 111646 3666
rect 115490 3614 115502 3666
rect 115554 3614 115566 3666
rect 73166 3602 73218 3614
rect 88510 3602 88562 3614
rect 94782 3602 94834 3614
rect 117406 3602 117458 3614
rect 2830 3554 2882 3566
rect 5954 3502 5966 3554
rect 6018 3502 6030 3554
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 10658 3502 10670 3554
rect 10722 3502 10734 3554
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 36306 3502 36318 3554
rect 36370 3502 36382 3554
rect 48850 3502 48862 3554
rect 48914 3502 48926 3554
rect 51650 3502 51662 3554
rect 51714 3502 51726 3554
rect 64978 3502 64990 3554
rect 65042 3502 65054 3554
rect 77522 3502 77534 3554
rect 77586 3502 77598 3554
rect 80882 3502 80894 3554
rect 80946 3502 80958 3554
rect 89954 3502 89966 3554
rect 90018 3502 90030 3554
rect 99810 3502 99822 3554
rect 99874 3502 99886 3554
rect 102610 3502 102622 3554
rect 102674 3502 102686 3554
rect 103842 3502 103854 3554
rect 103906 3502 103918 3554
rect 2830 3490 2882 3502
rect 2046 3442 2098 3454
rect 14590 3442 14642 3454
rect 24670 3442 24722 3454
rect 29374 3442 29426 3454
rect 41470 3442 41522 3454
rect 44270 3442 44322 3454
rect 53118 3442 53170 3454
rect 56590 3442 56642 3454
rect 3826 3390 3838 3442
rect 3890 3390 3902 3442
rect 9762 3390 9774 3442
rect 9826 3390 9838 3442
rect 15138 3390 15150 3442
rect 15202 3390 15214 3442
rect 19618 3390 19630 3442
rect 19682 3390 19694 3442
rect 21522 3390 21534 3442
rect 21586 3390 21598 3442
rect 25442 3390 25454 3442
rect 25506 3390 25518 3442
rect 29922 3390 29934 3442
rect 29986 3390 29998 3442
rect 37986 3390 37998 3442
rect 38050 3390 38062 3442
rect 42018 3390 42030 3442
rect 42082 3390 42094 3442
rect 45378 3390 45390 3442
rect 45442 3390 45454 3442
rect 50754 3390 50766 3442
rect 50818 3390 50830 3442
rect 55794 3390 55806 3442
rect 55858 3390 55870 3442
rect 2046 3378 2098 3390
rect 14590 3378 14642 3390
rect 24670 3378 24722 3390
rect 29374 3378 29426 3390
rect 41470 3378 41522 3390
rect 44270 3378 44322 3390
rect 53118 3378 53170 3390
rect 56590 3378 56642 3390
rect 57598 3442 57650 3454
rect 69022 3442 69074 3454
rect 83470 3442 83522 3454
rect 91310 3442 91362 3454
rect 95902 3442 95954 3454
rect 110910 3442 110962 3454
rect 114158 3442 114210 3454
rect 58146 3390 58158 3442
rect 58210 3390 58222 3442
rect 62738 3390 62750 3442
rect 62802 3390 62814 3442
rect 70466 3390 70478 3442
rect 70530 3390 70542 3442
rect 75058 3390 75070 3442
rect 75122 3390 75134 3442
rect 85138 3390 85150 3442
rect 85202 3390 85214 3442
rect 89058 3390 89070 3442
rect 89122 3390 89134 3442
rect 92978 3390 92990 3442
rect 93042 3390 93054 3442
rect 97346 3390 97358 3442
rect 97410 3390 97422 3442
rect 101714 3390 101726 3442
rect 101778 3390 101790 3442
rect 112578 3390 112590 3442
rect 112642 3390 112654 3442
rect 57598 3378 57650 3390
rect 69022 3378 69074 3390
rect 83470 3378 83522 3390
rect 91310 3378 91362 3390
rect 95902 3378 95954 3390
rect 110910 3378 110962 3390
rect 114158 3378 114210 3390
rect 114494 3442 114546 3454
rect 116498 3390 116510 3442
rect 116562 3390 116574 3442
rect 114494 3378 114546 3390
rect 2494 3330 2546 3342
rect 2494 3266 2546 3278
rect 27694 3330 27746 3342
rect 27694 3266 27746 3278
rect 28478 3330 28530 3342
rect 28478 3266 28530 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 76302 3330 76354 3342
rect 76302 3266 76354 3278
rect 80222 3330 80274 3342
rect 80222 3266 80274 3278
rect 105534 3330 105586 3342
rect 105534 3266 105586 3278
rect 109118 3330 109170 3342
rect 109118 3266 109170 3278
rect 109790 3330 109842 3342
rect 109790 3266 109842 3278
rect 118078 3330 118130 3342
rect 118078 3266 118130 3278
rect 1344 3162 118608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 118608 3162
rect 1344 3076 118608 3110
rect 104290 1710 104302 1762
rect 104354 1759 104366 1762
rect 105522 1759 105534 1762
rect 104354 1713 105534 1759
rect 104354 1710 104366 1713
rect 105522 1710 105534 1713
rect 105586 1710 105598 1762
<< via1 >>
rect 1710 117070 1762 117122
rect 1934 117070 1986 117122
rect 39790 117070 39842 117122
rect 41134 117070 41186 117122
rect 63982 116958 64034 117010
rect 65214 116958 65266 117010
rect 67230 116958 67282 117010
rect 68462 116958 68514 117010
rect 4478 116790 4530 116842
rect 4582 116790 4634 116842
rect 4686 116790 4738 116842
rect 35198 116790 35250 116842
rect 35302 116790 35354 116842
rect 35406 116790 35458 116842
rect 65918 116790 65970 116842
rect 66022 116790 66074 116842
rect 66126 116790 66178 116842
rect 96638 116790 96690 116842
rect 96742 116790 96794 116842
rect 96846 116790 96898 116842
rect 3278 116510 3330 116562
rect 5854 116510 5906 116562
rect 7534 116510 7586 116562
rect 9886 116510 9938 116562
rect 11790 116510 11842 116562
rect 12798 116510 12850 116562
rect 16718 116510 16770 116562
rect 21982 116510 22034 116562
rect 23886 116510 23938 116562
rect 26014 116510 26066 116562
rect 32174 116510 32226 116562
rect 36318 116510 36370 116562
rect 36990 116510 37042 116562
rect 37438 116510 37490 116562
rect 38110 116510 38162 116562
rect 39790 116510 39842 116562
rect 45054 116510 45106 116562
rect 48078 116510 48130 116562
rect 49534 116510 49586 116562
rect 51214 116510 51266 116562
rect 54014 116510 54066 116562
rect 56030 116510 56082 116562
rect 58158 116510 58210 116562
rect 59950 116510 60002 116562
rect 60958 116510 61010 116562
rect 65214 116510 65266 116562
rect 66446 116510 66498 116562
rect 69134 116510 69186 116562
rect 70590 116510 70642 116562
rect 72494 116510 72546 116562
rect 76974 116510 77026 116562
rect 78990 116510 79042 116562
rect 81118 116510 81170 116562
rect 81566 116510 81618 116562
rect 84814 116510 84866 116562
rect 86606 116510 86658 116562
rect 89070 116510 89122 116562
rect 92654 116510 92706 116562
rect 95118 116510 95170 116562
rect 95902 116510 95954 116562
rect 99150 116510 99202 116562
rect 99822 116510 99874 116562
rect 106878 116510 106930 116562
rect 107662 116510 107714 116562
rect 110910 116510 110962 116562
rect 111806 116510 111858 116562
rect 114830 116510 114882 116562
rect 115726 116510 115778 116562
rect 4062 116398 4114 116450
rect 17390 116398 17442 116450
rect 25342 116398 25394 116450
rect 53342 116398 53394 116450
rect 64542 116398 64594 116450
rect 67566 116398 67618 116450
rect 68462 116398 68514 116450
rect 71374 116398 71426 116450
rect 76302 116398 76354 116450
rect 78206 116398 78258 116450
rect 84142 116398 84194 116450
rect 85934 116398 85986 116450
rect 88286 116398 88338 116450
rect 91982 116398 92034 116450
rect 1934 116286 1986 116338
rect 6414 116286 6466 116338
rect 10446 116286 10498 116338
rect 15710 116286 15762 116338
rect 19070 116286 19122 116338
rect 22542 116286 22594 116338
rect 31390 116286 31442 116338
rect 33070 116286 33122 116338
rect 35198 116286 35250 116338
rect 38670 116286 38722 116338
rect 41134 116286 41186 116338
rect 44046 116286 44098 116338
rect 46958 116286 47010 116338
rect 48750 116286 48802 116338
rect 50094 116286 50146 116338
rect 56814 116286 56866 116338
rect 61742 116286 61794 116338
rect 74398 116286 74450 116338
rect 82574 116286 82626 116338
rect 94334 116286 94386 116338
rect 96910 116286 96962 116338
rect 97918 116286 97970 116338
rect 100830 116286 100882 116338
rect 108670 116286 108722 116338
rect 112814 116286 112866 116338
rect 116510 116286 116562 116338
rect 3838 116174 3890 116226
rect 4734 116174 4786 116226
rect 43598 116174 43650 116226
rect 52782 116174 52834 116226
rect 75518 116174 75570 116226
rect 91198 116174 91250 116226
rect 117518 116174 117570 116226
rect 19838 116006 19890 116058
rect 19942 116006 19994 116058
rect 20046 116006 20098 116058
rect 50558 116006 50610 116058
rect 50662 116006 50714 116058
rect 50766 116006 50818 116058
rect 81278 116006 81330 116058
rect 81382 116006 81434 116058
rect 81486 116006 81538 116058
rect 111998 116006 112050 116058
rect 112102 116006 112154 116058
rect 112206 116006 112258 116058
rect 5742 115838 5794 115890
rect 22766 115838 22818 115890
rect 23550 115838 23602 115890
rect 24110 115838 24162 115890
rect 28702 115838 28754 115890
rect 40798 115838 40850 115890
rect 41918 115838 41970 115890
rect 51326 115838 51378 115890
rect 67230 115838 67282 115890
rect 68686 115838 68738 115890
rect 69582 115838 69634 115890
rect 81790 115838 81842 115890
rect 85262 115838 85314 115890
rect 108670 115838 108722 115890
rect 1934 115726 1986 115778
rect 3726 115726 3778 115778
rect 10670 115726 10722 115778
rect 13134 115726 13186 115778
rect 29262 115726 29314 115778
rect 35310 115726 35362 115778
rect 37326 115726 37378 115778
rect 43598 115726 43650 115778
rect 45390 115726 45442 115778
rect 62862 115726 62914 115778
rect 72606 115726 72658 115778
rect 78990 115726 79042 115778
rect 83246 115726 83298 115778
rect 110126 115726 110178 115778
rect 111246 115726 111298 115778
rect 117854 115726 117906 115778
rect 3054 115614 3106 115666
rect 4622 115614 4674 115666
rect 10334 115614 10386 115666
rect 11230 115614 11282 115666
rect 23326 115614 23378 115666
rect 32846 115614 32898 115666
rect 36430 115614 36482 115666
rect 47294 115614 47346 115666
rect 56478 115614 56530 115666
rect 57822 115614 57874 115666
rect 59390 115614 59442 115666
rect 63982 115614 64034 115666
rect 67006 115614 67058 115666
rect 69022 115614 69074 115666
rect 71710 115614 71762 115666
rect 72382 115614 72434 115666
rect 73502 115614 73554 115666
rect 76862 115614 76914 115666
rect 80110 115614 80162 115666
rect 86270 115614 86322 115666
rect 87950 115614 88002 115666
rect 101054 115614 101106 115666
rect 112366 115614 112418 115666
rect 116174 115614 116226 115666
rect 116958 115614 117010 115666
rect 5294 115502 5346 115554
rect 9774 115502 9826 115554
rect 11902 115502 11954 115554
rect 14254 115502 14306 115554
rect 24670 115502 24722 115554
rect 30382 115502 30434 115554
rect 32062 115502 32114 115554
rect 33630 115502 33682 115554
rect 38670 115502 38722 115554
rect 44494 115502 44546 115554
rect 46510 115502 46562 115554
rect 47966 115502 48018 115554
rect 55694 115502 55746 115554
rect 58270 115502 58322 115554
rect 60062 115502 60114 115554
rect 64430 115502 64482 115554
rect 66334 115502 66386 115554
rect 70142 115502 70194 115554
rect 71262 115502 71314 115554
rect 74174 115502 74226 115554
rect 76414 115502 76466 115554
rect 77534 115502 77586 115554
rect 80558 115502 80610 115554
rect 82238 115502 82290 115554
rect 84142 115502 84194 115554
rect 85822 115502 85874 115554
rect 86942 115502 86994 115554
rect 100494 115502 100546 115554
rect 101726 115502 101778 115554
rect 109118 115502 109170 115554
rect 115502 115502 115554 115554
rect 4478 115222 4530 115274
rect 4582 115222 4634 115274
rect 4686 115222 4738 115274
rect 35198 115222 35250 115274
rect 35302 115222 35354 115274
rect 35406 115222 35458 115274
rect 65918 115222 65970 115274
rect 66022 115222 66074 115274
rect 66126 115222 66178 115274
rect 96638 115222 96690 115274
rect 96742 115222 96794 115274
rect 96846 115222 96898 115274
rect 2046 114942 2098 114994
rect 4398 114942 4450 114994
rect 11342 114942 11394 114994
rect 12350 114942 12402 114994
rect 33966 114942 34018 114994
rect 36654 114942 36706 114994
rect 45390 114942 45442 114994
rect 46958 114942 47010 114994
rect 59166 114942 59218 114994
rect 62974 114942 63026 114994
rect 72158 114942 72210 114994
rect 77870 114942 77922 114994
rect 115838 114942 115890 114994
rect 3054 114830 3106 114882
rect 3614 114830 3666 114882
rect 11902 114830 11954 114882
rect 34862 114830 34914 114882
rect 63646 114830 63698 114882
rect 64430 114830 64482 114882
rect 110798 114830 110850 114882
rect 114382 114830 114434 114882
rect 115166 114830 115218 114882
rect 117294 114830 117346 114882
rect 3950 114718 4002 114770
rect 56926 114718 56978 114770
rect 57486 114718 57538 114770
rect 57822 114718 57874 114770
rect 63870 114718 63922 114770
rect 64766 114718 64818 114770
rect 86942 114718 86994 114770
rect 117070 114718 117122 114770
rect 23774 114606 23826 114658
rect 35534 114606 35586 114658
rect 56478 114606 56530 114658
rect 19838 114438 19890 114490
rect 19942 114438 19994 114490
rect 20046 114438 20098 114490
rect 50558 114438 50610 114490
rect 50662 114438 50714 114490
rect 50766 114438 50818 114490
rect 81278 114438 81330 114490
rect 81382 114438 81434 114490
rect 81486 114438 81538 114490
rect 111998 114438 112050 114490
rect 112102 114438 112154 114490
rect 112206 114438 112258 114490
rect 64094 114270 64146 114322
rect 117070 114270 117122 114322
rect 1934 114158 1986 114210
rect 3726 114046 3778 114098
rect 116174 114046 116226 114098
rect 3278 113934 3330 113986
rect 115502 113934 115554 113986
rect 116174 113934 116226 113986
rect 116734 113934 116786 113986
rect 116734 113822 116786 113874
rect 4478 113654 4530 113706
rect 4582 113654 4634 113706
rect 4686 113654 4738 113706
rect 35198 113654 35250 113706
rect 35302 113654 35354 113706
rect 35406 113654 35458 113706
rect 65918 113654 65970 113706
rect 66022 113654 66074 113706
rect 66126 113654 66178 113706
rect 96638 113654 96690 113706
rect 96742 113654 96794 113706
rect 96846 113654 96898 113706
rect 1822 113374 1874 113426
rect 2830 113150 2882 113202
rect 2494 113038 2546 113090
rect 3278 113038 3330 113090
rect 19838 112870 19890 112922
rect 19942 112870 19994 112922
rect 20046 112870 20098 112922
rect 50558 112870 50610 112922
rect 50662 112870 50714 112922
rect 50766 112870 50818 112922
rect 81278 112870 81330 112922
rect 81382 112870 81434 112922
rect 81486 112870 81538 112922
rect 111998 112870 112050 112922
rect 112102 112870 112154 112922
rect 112206 112870 112258 112922
rect 118078 112590 118130 112642
rect 2830 112478 2882 112530
rect 1934 112366 1986 112418
rect 4478 112086 4530 112138
rect 4582 112086 4634 112138
rect 4686 112086 4738 112138
rect 35198 112086 35250 112138
rect 35302 112086 35354 112138
rect 35406 112086 35458 112138
rect 65918 112086 65970 112138
rect 66022 112086 66074 112138
rect 66126 112086 66178 112138
rect 96638 112086 96690 112138
rect 96742 112086 96794 112138
rect 96846 112086 96898 112138
rect 3278 111806 3330 111858
rect 1934 111582 1986 111634
rect 118078 111470 118130 111522
rect 19838 111302 19890 111354
rect 19942 111302 19994 111354
rect 20046 111302 20098 111354
rect 50558 111302 50610 111354
rect 50662 111302 50714 111354
rect 50766 111302 50818 111354
rect 81278 111302 81330 111354
rect 81382 111302 81434 111354
rect 81486 111302 81538 111354
rect 111998 111302 112050 111354
rect 112102 111302 112154 111354
rect 112206 111302 112258 111354
rect 1710 111022 1762 111074
rect 115166 110910 115218 110962
rect 115838 110798 115890 110850
rect 116622 110798 116674 110850
rect 4478 110518 4530 110570
rect 4582 110518 4634 110570
rect 4686 110518 4738 110570
rect 35198 110518 35250 110570
rect 35302 110518 35354 110570
rect 35406 110518 35458 110570
rect 65918 110518 65970 110570
rect 66022 110518 66074 110570
rect 66126 110518 66178 110570
rect 96638 110518 96690 110570
rect 96742 110518 96794 110570
rect 96846 110518 96898 110570
rect 1822 109902 1874 109954
rect 19838 109734 19890 109786
rect 19942 109734 19994 109786
rect 20046 109734 20098 109786
rect 50558 109734 50610 109786
rect 50662 109734 50714 109786
rect 50766 109734 50818 109786
rect 81278 109734 81330 109786
rect 81382 109734 81434 109786
rect 81486 109734 81538 109786
rect 111998 109734 112050 109786
rect 112102 109734 112154 109786
rect 112206 109734 112258 109786
rect 116286 109454 116338 109506
rect 114942 109230 114994 109282
rect 116846 109230 116898 109282
rect 4478 108950 4530 109002
rect 4582 108950 4634 109002
rect 4686 108950 4738 109002
rect 35198 108950 35250 109002
rect 35302 108950 35354 109002
rect 35406 108950 35458 109002
rect 65918 108950 65970 109002
rect 66022 108950 66074 109002
rect 66126 108950 66178 109002
rect 96638 108950 96690 109002
rect 96742 108950 96794 109002
rect 96846 108950 96898 109002
rect 19838 108166 19890 108218
rect 19942 108166 19994 108218
rect 20046 108166 20098 108218
rect 50558 108166 50610 108218
rect 50662 108166 50714 108218
rect 50766 108166 50818 108218
rect 81278 108166 81330 108218
rect 81382 108166 81434 108218
rect 81486 108166 81538 108218
rect 111998 108166 112050 108218
rect 112102 108166 112154 108218
rect 112206 108166 112258 108218
rect 1822 107886 1874 107938
rect 116286 107886 116338 107938
rect 114942 107662 114994 107714
rect 116846 107662 116898 107714
rect 4478 107382 4530 107434
rect 4582 107382 4634 107434
rect 4686 107382 4738 107434
rect 35198 107382 35250 107434
rect 35302 107382 35354 107434
rect 35406 107382 35458 107434
rect 65918 107382 65970 107434
rect 66022 107382 66074 107434
rect 66126 107382 66178 107434
rect 96638 107382 96690 107434
rect 96742 107382 96794 107434
rect 96846 107382 96898 107434
rect 118078 106766 118130 106818
rect 19838 106598 19890 106650
rect 19942 106598 19994 106650
rect 20046 106598 20098 106650
rect 50558 106598 50610 106650
rect 50662 106598 50714 106650
rect 50766 106598 50818 106650
rect 81278 106598 81330 106650
rect 81382 106598 81434 106650
rect 81486 106598 81538 106650
rect 111998 106598 112050 106650
rect 112102 106598 112154 106650
rect 112206 106598 112258 106650
rect 114494 106206 114546 106258
rect 114942 106206 114994 106258
rect 115838 106094 115890 106146
rect 4478 105814 4530 105866
rect 4582 105814 4634 105866
rect 4686 105814 4738 105866
rect 35198 105814 35250 105866
rect 35302 105814 35354 105866
rect 35406 105814 35458 105866
rect 65918 105814 65970 105866
rect 66022 105814 66074 105866
rect 66126 105814 66178 105866
rect 96638 105814 96690 105866
rect 96742 105814 96794 105866
rect 96846 105814 96898 105866
rect 19838 105030 19890 105082
rect 19942 105030 19994 105082
rect 20046 105030 20098 105082
rect 50558 105030 50610 105082
rect 50662 105030 50714 105082
rect 50766 105030 50818 105082
rect 81278 105030 81330 105082
rect 81382 105030 81434 105082
rect 81486 105030 81538 105082
rect 111998 105030 112050 105082
rect 112102 105030 112154 105082
rect 112206 105030 112258 105082
rect 116286 104750 116338 104802
rect 3054 104638 3106 104690
rect 1934 104526 1986 104578
rect 3614 104526 3666 104578
rect 114942 104526 114994 104578
rect 116846 104526 116898 104578
rect 4478 104246 4530 104298
rect 4582 104246 4634 104298
rect 4686 104246 4738 104298
rect 35198 104246 35250 104298
rect 35302 104246 35354 104298
rect 35406 104246 35458 104298
rect 65918 104246 65970 104298
rect 66022 104246 66074 104298
rect 66126 104246 66178 104298
rect 96638 104246 96690 104298
rect 96742 104246 96794 104298
rect 96846 104246 96898 104298
rect 19838 103462 19890 103514
rect 19942 103462 19994 103514
rect 20046 103462 20098 103514
rect 50558 103462 50610 103514
rect 50662 103462 50714 103514
rect 50766 103462 50818 103514
rect 81278 103462 81330 103514
rect 81382 103462 81434 103514
rect 81486 103462 81538 103514
rect 111998 103462 112050 103514
rect 112102 103462 112154 103514
rect 112206 103462 112258 103514
rect 44830 103182 44882 103234
rect 3054 103070 3106 103122
rect 45166 103070 45218 103122
rect 1934 102958 1986 103010
rect 3614 102958 3666 103010
rect 45614 102958 45666 103010
rect 4478 102678 4530 102730
rect 4582 102678 4634 102730
rect 4686 102678 4738 102730
rect 35198 102678 35250 102730
rect 35302 102678 35354 102730
rect 35406 102678 35458 102730
rect 65918 102678 65970 102730
rect 66022 102678 66074 102730
rect 66126 102678 66178 102730
rect 96638 102678 96690 102730
rect 96742 102678 96794 102730
rect 96846 102678 96898 102730
rect 3166 102398 3218 102450
rect 114830 102398 114882 102450
rect 2270 102174 2322 102226
rect 116062 102174 116114 102226
rect 117070 102062 117122 102114
rect 19838 101894 19890 101946
rect 19942 101894 19994 101946
rect 20046 101894 20098 101946
rect 50558 101894 50610 101946
rect 50662 101894 50714 101946
rect 50766 101894 50818 101946
rect 81278 101894 81330 101946
rect 81382 101894 81434 101946
rect 81486 101894 81538 101946
rect 111998 101894 112050 101946
rect 112102 101894 112154 101946
rect 112206 101894 112258 101946
rect 1822 101614 1874 101666
rect 2382 101614 2434 101666
rect 118078 101614 118130 101666
rect 4478 101110 4530 101162
rect 4582 101110 4634 101162
rect 4686 101110 4738 101162
rect 35198 101110 35250 101162
rect 35302 101110 35354 101162
rect 35406 101110 35458 101162
rect 65918 101110 65970 101162
rect 66022 101110 66074 101162
rect 66126 101110 66178 101162
rect 96638 101110 96690 101162
rect 96742 101110 96794 101162
rect 96846 101110 96898 101162
rect 19838 100326 19890 100378
rect 19942 100326 19994 100378
rect 20046 100326 20098 100378
rect 50558 100326 50610 100378
rect 50662 100326 50714 100378
rect 50766 100326 50818 100378
rect 81278 100326 81330 100378
rect 81382 100326 81434 100378
rect 81486 100326 81538 100378
rect 111998 100326 112050 100378
rect 112102 100326 112154 100378
rect 112206 100326 112258 100378
rect 1934 100046 1986 100098
rect 114494 99934 114546 99986
rect 114942 99934 114994 99986
rect 3278 99822 3330 99874
rect 115838 99822 115890 99874
rect 4478 99542 4530 99594
rect 4582 99542 4634 99594
rect 4686 99542 4738 99594
rect 35198 99542 35250 99594
rect 35302 99542 35354 99594
rect 35406 99542 35458 99594
rect 65918 99542 65970 99594
rect 66022 99542 66074 99594
rect 66126 99542 66178 99594
rect 96638 99542 96690 99594
rect 96742 99542 96794 99594
rect 96846 99542 96898 99594
rect 38558 99374 38610 99426
rect 1822 99262 1874 99314
rect 37886 99262 37938 99314
rect 38334 99262 38386 99314
rect 39454 99262 39506 99314
rect 2606 99150 2658 99202
rect 38894 99150 38946 99202
rect 2830 98926 2882 98978
rect 3278 98926 3330 98978
rect 19838 98758 19890 98810
rect 19942 98758 19994 98810
rect 20046 98758 20098 98810
rect 50558 98758 50610 98810
rect 50662 98758 50714 98810
rect 50766 98758 50818 98810
rect 81278 98758 81330 98810
rect 81382 98758 81434 98810
rect 81486 98758 81538 98810
rect 111998 98758 112050 98810
rect 112102 98758 112154 98810
rect 112206 98758 112258 98810
rect 2830 98366 2882 98418
rect 1934 98254 1986 98306
rect 4478 97974 4530 98026
rect 4582 97974 4634 98026
rect 4686 97974 4738 98026
rect 35198 97974 35250 98026
rect 35302 97974 35354 98026
rect 35406 97974 35458 98026
rect 65918 97974 65970 98026
rect 66022 97974 66074 98026
rect 66126 97974 66178 98026
rect 96638 97974 96690 98026
rect 96742 97974 96794 98026
rect 96846 97974 96898 98026
rect 3278 97694 3330 97746
rect 1934 97470 1986 97522
rect 19838 97190 19890 97242
rect 19942 97190 19994 97242
rect 20046 97190 20098 97242
rect 50558 97190 50610 97242
rect 50662 97190 50714 97242
rect 50766 97190 50818 97242
rect 81278 97190 81330 97242
rect 81382 97190 81434 97242
rect 81486 97190 81538 97242
rect 111998 97190 112050 97242
rect 112102 97190 112154 97242
rect 112206 97190 112258 97242
rect 1710 96910 1762 96962
rect 118078 96910 118130 96962
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 65918 96406 65970 96458
rect 66022 96406 66074 96458
rect 66126 96406 66178 96458
rect 96638 96406 96690 96458
rect 96742 96406 96794 96458
rect 96846 96406 96898 96458
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 50558 95622 50610 95674
rect 50662 95622 50714 95674
rect 50766 95622 50818 95674
rect 81278 95622 81330 95674
rect 81382 95622 81434 95674
rect 81486 95622 81538 95674
rect 111998 95622 112050 95674
rect 112102 95622 112154 95674
rect 112206 95622 112258 95674
rect 2830 95230 2882 95282
rect 114942 95230 114994 95282
rect 1934 95118 1986 95170
rect 114494 95118 114546 95170
rect 115838 95118 115890 95170
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 65918 94838 65970 94890
rect 66022 94838 66074 94890
rect 66126 94838 66178 94890
rect 96638 94838 96690 94890
rect 96742 94838 96794 94890
rect 96846 94838 96898 94890
rect 3278 94558 3330 94610
rect 114830 94558 114882 94610
rect 2830 94446 2882 94498
rect 2494 94334 2546 94386
rect 71262 94334 71314 94386
rect 71822 94334 71874 94386
rect 116062 94334 116114 94386
rect 72158 94222 72210 94274
rect 117070 94222 117122 94274
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 50558 94054 50610 94106
rect 50662 94054 50714 94106
rect 50766 94054 50818 94106
rect 81278 94054 81330 94106
rect 81382 94054 81434 94106
rect 81486 94054 81538 94106
rect 111998 94054 112050 94106
rect 112102 94054 112154 94106
rect 112206 94054 112258 94106
rect 48302 93774 48354 93826
rect 3054 93662 3106 93714
rect 48638 93662 48690 93714
rect 1934 93550 1986 93602
rect 3614 93550 3666 93602
rect 49422 93550 49474 93602
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 65918 93270 65970 93322
rect 66022 93270 66074 93322
rect 66126 93270 66178 93322
rect 96638 93270 96690 93322
rect 96742 93270 96794 93322
rect 96846 93270 96898 93322
rect 3278 92990 3330 93042
rect 115838 92990 115890 93042
rect 114382 92878 114434 92930
rect 114942 92878 114994 92930
rect 1934 92766 1986 92818
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 50558 92486 50610 92538
rect 50662 92486 50714 92538
rect 50766 92486 50818 92538
rect 81278 92486 81330 92538
rect 81382 92486 81434 92538
rect 81486 92486 81538 92538
rect 111998 92486 112050 92538
rect 112102 92486 112154 92538
rect 112206 92486 112258 92538
rect 1822 92318 1874 92370
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 65918 91702 65970 91754
rect 66022 91702 66074 91754
rect 66126 91702 66178 91754
rect 96638 91702 96690 91754
rect 96742 91702 96794 91754
rect 96846 91702 96898 91754
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 50558 90918 50610 90970
rect 50662 90918 50714 90970
rect 50766 90918 50818 90970
rect 81278 90918 81330 90970
rect 81382 90918 81434 90970
rect 81486 90918 81538 90970
rect 111998 90918 112050 90970
rect 112102 90918 112154 90970
rect 112206 90918 112258 90970
rect 2830 90526 2882 90578
rect 1934 90414 1986 90466
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 65918 90134 65970 90186
rect 66022 90134 66074 90186
rect 66126 90134 66178 90186
rect 96638 90134 96690 90186
rect 96742 90134 96794 90186
rect 96846 90134 96898 90186
rect 3054 89966 3106 90018
rect 3278 89966 3330 90018
rect 3278 89854 3330 89906
rect 115390 89854 115442 89906
rect 2830 89742 2882 89794
rect 115950 89742 116002 89794
rect 2494 89630 2546 89682
rect 58830 89630 58882 89682
rect 59166 89630 59218 89682
rect 116958 89630 117010 89682
rect 59726 89518 59778 89570
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 50558 89350 50610 89402
rect 50662 89350 50714 89402
rect 50766 89350 50818 89402
rect 81278 89350 81330 89402
rect 81382 89350 81434 89402
rect 81486 89350 81538 89402
rect 111998 89350 112050 89402
rect 112102 89350 112154 89402
rect 112206 89350 112258 89402
rect 3054 88958 3106 89010
rect 3502 88958 3554 89010
rect 1934 88846 1986 88898
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 65918 88566 65970 88618
rect 66022 88566 66074 88618
rect 66126 88566 66178 88618
rect 96638 88566 96690 88618
rect 96742 88566 96794 88618
rect 96846 88566 96898 88618
rect 3278 88286 3330 88338
rect 1934 88062 1986 88114
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 50558 87782 50610 87834
rect 50662 87782 50714 87834
rect 50766 87782 50818 87834
rect 81278 87782 81330 87834
rect 81382 87782 81434 87834
rect 81486 87782 81538 87834
rect 111998 87782 112050 87834
rect 112102 87782 112154 87834
rect 112206 87782 112258 87834
rect 1822 87614 1874 87666
rect 116286 87502 116338 87554
rect 116846 87390 116898 87442
rect 114942 87278 114994 87330
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 65918 86998 65970 87050
rect 66022 86998 66074 87050
rect 66126 86998 66178 87050
rect 96638 86998 96690 87050
rect 96742 86998 96794 87050
rect 96846 86998 96898 87050
rect 115838 86718 115890 86770
rect 114382 86606 114434 86658
rect 114942 86606 114994 86658
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 50558 86214 50610 86266
rect 50662 86214 50714 86266
rect 50766 86214 50818 86266
rect 81278 86214 81330 86266
rect 81382 86214 81434 86266
rect 81486 86214 81538 86266
rect 111998 86214 112050 86266
rect 112102 86214 112154 86266
rect 112206 86214 112258 86266
rect 1822 85934 1874 85986
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 65918 85430 65970 85482
rect 66022 85430 66074 85482
rect 66126 85430 66178 85482
rect 96638 85430 96690 85482
rect 96742 85430 96794 85482
rect 96846 85430 96898 85482
rect 115838 85150 115890 85202
rect 114494 85038 114546 85090
rect 114942 85038 114994 85090
rect 76190 84926 76242 84978
rect 75630 84814 75682 84866
rect 76526 84814 76578 84866
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 50558 84646 50610 84698
rect 50662 84646 50714 84698
rect 50766 84646 50818 84698
rect 81278 84646 81330 84698
rect 81382 84646 81434 84698
rect 81486 84646 81538 84698
rect 111998 84646 112050 84698
rect 112102 84646 112154 84698
rect 112206 84646 112258 84698
rect 1822 84366 1874 84418
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 65918 83862 65970 83914
rect 66022 83862 66074 83914
rect 66126 83862 66178 83914
rect 96638 83862 96690 83914
rect 96742 83862 96794 83914
rect 96846 83862 96898 83914
rect 115390 83582 115442 83634
rect 116174 83470 116226 83522
rect 117294 83470 117346 83522
rect 117070 83358 117122 83410
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 50558 83078 50610 83130
rect 50662 83078 50714 83130
rect 50766 83078 50818 83130
rect 81278 83078 81330 83130
rect 81382 83078 81434 83130
rect 81486 83078 81538 83130
rect 111998 83078 112050 83130
rect 112102 83078 112154 83130
rect 112206 83078 112258 83130
rect 116734 82910 116786 82962
rect 118078 82798 118130 82850
rect 2830 82686 2882 82738
rect 1934 82574 1986 82626
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 65918 82294 65970 82346
rect 66022 82294 66074 82346
rect 66126 82294 66178 82346
rect 96638 82294 96690 82346
rect 96742 82294 96794 82346
rect 96846 82294 96898 82346
rect 3054 82126 3106 82178
rect 3278 82126 3330 82178
rect 3278 82014 3330 82066
rect 2830 81902 2882 81954
rect 2494 81790 2546 81842
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 50558 81510 50610 81562
rect 50662 81510 50714 81562
rect 50766 81510 50818 81562
rect 81278 81510 81330 81562
rect 81382 81510 81434 81562
rect 81486 81510 81538 81562
rect 111998 81510 112050 81562
rect 112102 81510 112154 81562
rect 112206 81510 112258 81562
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 65918 80726 65970 80778
rect 66022 80726 66074 80778
rect 66126 80726 66178 80778
rect 96638 80726 96690 80778
rect 96742 80726 96794 80778
rect 96846 80726 96898 80778
rect 2830 80334 2882 80386
rect 1934 80222 1986 80274
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 50558 79942 50610 79994
rect 50662 79942 50714 79994
rect 50766 79942 50818 79994
rect 81278 79942 81330 79994
rect 81382 79942 81434 79994
rect 81486 79942 81538 79994
rect 111998 79942 112050 79994
rect 112102 79942 112154 79994
rect 112206 79942 112258 79994
rect 2494 79774 2546 79826
rect 3278 79774 3330 79826
rect 117966 79774 118018 79826
rect 117294 79662 117346 79714
rect 2830 79550 2882 79602
rect 3054 79326 3106 79378
rect 3278 79326 3330 79378
rect 114830 79326 114882 79378
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 65918 79158 65970 79210
rect 66022 79158 66074 79210
rect 66126 79158 66178 79210
rect 96638 79158 96690 79210
rect 96742 79158 96794 79210
rect 96846 79158 96898 79210
rect 3054 78766 3106 78818
rect 1934 78654 1986 78706
rect 3502 78542 3554 78594
rect 118078 78542 118130 78594
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 50558 78374 50610 78426
rect 50662 78374 50714 78426
rect 50766 78374 50818 78426
rect 81278 78374 81330 78426
rect 81382 78374 81434 78426
rect 81486 78374 81538 78426
rect 111998 78374 112050 78426
rect 112102 78374 112154 78426
rect 112206 78374 112258 78426
rect 117966 78206 118018 78258
rect 117182 78094 117234 78146
rect 114830 77758 114882 77810
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 65918 77590 65970 77642
rect 66022 77590 66074 77642
rect 66126 77590 66178 77642
rect 96638 77590 96690 77642
rect 96742 77590 96794 77642
rect 96846 77590 96898 77642
rect 1822 76974 1874 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 81278 76806 81330 76858
rect 81382 76806 81434 76858
rect 81486 76806 81538 76858
rect 111998 76806 112050 76858
rect 112102 76806 112154 76858
rect 112206 76806 112258 76858
rect 1934 76526 1986 76578
rect 4398 76190 4450 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 96638 76022 96690 76074
rect 96742 76022 96794 76074
rect 96846 76022 96898 76074
rect 2830 75630 2882 75682
rect 114382 75630 114434 75682
rect 114942 75630 114994 75682
rect 1934 75518 1986 75570
rect 116062 75518 116114 75570
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 81278 75238 81330 75290
rect 81382 75238 81434 75290
rect 81486 75238 81538 75290
rect 111998 75238 112050 75290
rect 112102 75238 112154 75290
rect 112206 75238 112258 75290
rect 2494 75070 2546 75122
rect 3278 75070 3330 75122
rect 2830 74958 2882 75010
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 96638 74454 96690 74506
rect 96742 74454 96794 74506
rect 96846 74454 96898 74506
rect 114830 74174 114882 74226
rect 116174 73950 116226 74002
rect 117070 73950 117122 74002
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 81278 73670 81330 73722
rect 81382 73670 81434 73722
rect 81486 73670 81538 73722
rect 111998 73670 112050 73722
rect 112102 73670 112154 73722
rect 112206 73670 112258 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 96638 72886 96690 72938
rect 96742 72886 96794 72938
rect 96846 72886 96898 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 81278 72102 81330 72154
rect 81382 72102 81434 72154
rect 81486 72102 81538 72154
rect 111998 72102 112050 72154
rect 112102 72102 112154 72154
rect 112206 72102 112258 72154
rect 1934 71822 1986 71874
rect 3278 71598 3330 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 96638 71318 96690 71370
rect 96742 71318 96794 71370
rect 96846 71318 96898 71370
rect 1822 71038 1874 71090
rect 118078 70702 118130 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 81278 70534 81330 70586
rect 81382 70534 81434 70586
rect 81486 70534 81538 70586
rect 111998 70534 112050 70586
rect 112102 70534 112154 70586
rect 112206 70534 112258 70586
rect 3390 70366 3442 70418
rect 115502 70366 115554 70418
rect 115950 70366 116002 70418
rect 2494 70254 2546 70306
rect 2830 70254 2882 70306
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 96638 69750 96690 69802
rect 96742 69750 96794 69802
rect 96846 69750 96898 69802
rect 115838 69470 115890 69522
rect 2830 69358 2882 69410
rect 114382 69358 114434 69410
rect 114942 69358 114994 69410
rect 1934 69246 1986 69298
rect 55918 69134 55970 69186
rect 117070 69134 117122 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 81278 68966 81330 69018
rect 81382 68966 81434 69018
rect 81486 68966 81538 69018
rect 111998 68966 112050 69018
rect 112102 68966 112154 69018
rect 112206 68966 112258 69018
rect 46398 68798 46450 68850
rect 116398 68686 116450 68738
rect 116958 68686 117010 68738
rect 3054 68574 3106 68626
rect 46062 68574 46114 68626
rect 114494 68574 114546 68626
rect 1934 68462 1986 68514
rect 3614 68462 3666 68514
rect 46846 68462 46898 68514
rect 55246 68462 55298 68514
rect 55694 68462 55746 68514
rect 56142 68462 56194 68514
rect 56478 68462 56530 68514
rect 63086 68462 63138 68514
rect 63982 68462 64034 68514
rect 114046 68462 114098 68514
rect 115614 68462 115666 68514
rect 117182 68350 117234 68402
rect 117518 68350 117570 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 96638 68182 96690 68234
rect 96742 68182 96794 68234
rect 96846 68182 96898 68234
rect 57038 68014 57090 68066
rect 54910 67902 54962 67954
rect 56590 67902 56642 67954
rect 60622 67902 60674 67954
rect 63646 67902 63698 67954
rect 64094 67902 64146 67954
rect 115502 67902 115554 67954
rect 49310 67790 49362 67842
rect 55134 67790 55186 67842
rect 56702 67790 56754 67842
rect 61854 67790 61906 67842
rect 62638 67790 62690 67842
rect 74846 67790 74898 67842
rect 77534 67790 77586 67842
rect 116174 67790 116226 67842
rect 117406 67790 117458 67842
rect 55694 67678 55746 67730
rect 62526 67678 62578 67730
rect 63310 67678 63362 67730
rect 71710 67678 71762 67730
rect 77758 67678 77810 67730
rect 49646 67566 49698 67618
rect 57822 67566 57874 67618
rect 61518 67566 61570 67618
rect 63534 67566 63586 67618
rect 64542 67566 64594 67618
rect 72046 67566 72098 67618
rect 75070 67566 75122 67618
rect 78318 67566 78370 67618
rect 117070 67566 117122 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 81278 67398 81330 67450
rect 81382 67398 81434 67450
rect 81486 67398 81538 67450
rect 111998 67398 112050 67450
rect 112102 67398 112154 67450
rect 112206 67398 112258 67450
rect 56590 67230 56642 67282
rect 71374 67230 71426 67282
rect 82350 67230 82402 67282
rect 48638 67118 48690 67170
rect 50542 67118 50594 67170
rect 56254 67118 56306 67170
rect 56366 67118 56418 67170
rect 72270 67118 72322 67170
rect 74958 67118 75010 67170
rect 78430 67118 78482 67170
rect 117294 67118 117346 67170
rect 48414 67006 48466 67058
rect 49646 67006 49698 67058
rect 50766 67006 50818 67058
rect 52670 67006 52722 67058
rect 57598 67006 57650 67058
rect 61294 67006 61346 67058
rect 65326 67006 65378 67058
rect 72382 67006 72434 67058
rect 74286 67006 74338 67058
rect 77646 67006 77698 67058
rect 82014 67006 82066 67058
rect 117966 67006 118018 67058
rect 51326 66894 51378 66946
rect 53342 66894 53394 66946
rect 55582 66894 55634 66946
rect 58270 66894 58322 66946
rect 60510 66894 60562 66946
rect 61966 66894 62018 66946
rect 64094 66894 64146 66946
rect 64542 66894 64594 66946
rect 70254 66894 70306 66946
rect 70702 66894 70754 66946
rect 73278 66894 73330 66946
rect 77086 66894 77138 66946
rect 80558 66894 80610 66946
rect 81230 66894 81282 66946
rect 113934 66894 113986 66946
rect 114382 66894 114434 66946
rect 115166 66894 115218 66946
rect 49982 66782 50034 66834
rect 71710 66782 71762 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 96638 66614 96690 66666
rect 96742 66614 96794 66666
rect 96846 66614 96898 66666
rect 53678 66446 53730 66498
rect 74846 66446 74898 66498
rect 76302 66446 76354 66498
rect 76526 66446 76578 66498
rect 77870 66446 77922 66498
rect 3278 66334 3330 66386
rect 47294 66334 47346 66386
rect 49422 66334 49474 66386
rect 55470 66334 55522 66386
rect 55918 66334 55970 66386
rect 57262 66334 57314 66386
rect 58270 66334 58322 66386
rect 58942 66334 58994 66386
rect 59390 66334 59442 66386
rect 60622 66334 60674 66386
rect 63758 66334 63810 66386
rect 65886 66334 65938 66386
rect 72046 66334 72098 66386
rect 74174 66334 74226 66386
rect 76526 66334 76578 66386
rect 79550 66334 79602 66386
rect 45614 66222 45666 66274
rect 50206 66222 50258 66274
rect 54574 66222 54626 66274
rect 54798 66222 54850 66274
rect 54910 66222 54962 66274
rect 55246 66222 55298 66274
rect 56590 66222 56642 66274
rect 56702 66222 56754 66274
rect 57038 66222 57090 66274
rect 57598 66222 57650 66274
rect 58494 66222 58546 66274
rect 61518 66222 61570 66274
rect 62974 66222 63026 66274
rect 71374 66222 71426 66274
rect 75182 66222 75234 66274
rect 75630 66222 75682 66274
rect 78206 66222 78258 66274
rect 114158 66222 114210 66274
rect 115054 66222 115106 66274
rect 115390 66222 115442 66274
rect 117406 66222 117458 66274
rect 1934 66110 1986 66162
rect 52334 66110 52386 66162
rect 52670 66110 52722 66162
rect 54014 66110 54066 66162
rect 58158 66110 58210 66162
rect 61742 66110 61794 66162
rect 75966 66110 76018 66162
rect 77198 66110 77250 66162
rect 78430 66110 78482 66162
rect 78878 66110 78930 66162
rect 113486 66110 113538 66162
rect 115614 66110 115666 66162
rect 116062 66110 116114 66162
rect 117070 66110 117122 66162
rect 117854 66110 117906 66162
rect 45838 65998 45890 66050
rect 50654 65998 50706 66050
rect 51886 65998 51938 66050
rect 53790 65998 53842 66050
rect 55358 65998 55410 66050
rect 56478 65998 56530 66050
rect 57710 65998 57762 66050
rect 62190 65998 62242 66050
rect 66334 65998 66386 66050
rect 66782 65998 66834 66050
rect 67342 65998 67394 66050
rect 69246 65998 69298 66050
rect 81678 65998 81730 66050
rect 114382 65998 114434 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 81278 65830 81330 65882
rect 81382 65830 81434 65882
rect 81486 65830 81538 65882
rect 111998 65830 112050 65882
rect 112102 65830 112154 65882
rect 112206 65830 112258 65882
rect 1822 65662 1874 65714
rect 54686 65662 54738 65714
rect 55022 65662 55074 65714
rect 55582 65662 55634 65714
rect 63310 65662 63362 65714
rect 77422 65662 77474 65714
rect 113934 65662 113986 65714
rect 46734 65550 46786 65602
rect 58494 65550 58546 65602
rect 62302 65550 62354 65602
rect 115278 65550 115330 65602
rect 47518 65438 47570 65490
rect 47966 65438 48018 65490
rect 49534 65438 49586 65490
rect 49982 65438 50034 65490
rect 53342 65438 53394 65490
rect 61518 65438 61570 65490
rect 62414 65438 62466 65490
rect 62526 65438 62578 65490
rect 62974 65438 63026 65490
rect 64654 65438 64706 65490
rect 65662 65438 65714 65490
rect 69134 65438 69186 65490
rect 74622 65438 74674 65490
rect 114494 65438 114546 65490
rect 117854 65438 117906 65490
rect 44606 65326 44658 65378
rect 48750 65326 48802 65378
rect 53790 65326 53842 65378
rect 54238 65326 54290 65378
rect 55918 65326 55970 65378
rect 56142 65326 56194 65378
rect 56590 65326 56642 65378
rect 57486 65326 57538 65378
rect 58046 65326 58098 65378
rect 59838 65326 59890 65378
rect 60958 65326 61010 65378
rect 63198 65326 63250 65378
rect 63534 65326 63586 65378
rect 63870 65326 63922 65378
rect 66446 65326 66498 65378
rect 68574 65326 68626 65378
rect 69918 65326 69970 65378
rect 72046 65326 72098 65378
rect 74174 65326 74226 65378
rect 75070 65326 75122 65378
rect 117406 65326 117458 65378
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 96638 65046 96690 65098
rect 96742 65046 96794 65098
rect 96846 65046 96898 65098
rect 45614 64878 45666 64930
rect 62190 64878 62242 64930
rect 62526 64878 62578 64930
rect 44718 64766 44770 64818
rect 54910 64766 54962 64818
rect 57150 64766 57202 64818
rect 60174 64766 60226 64818
rect 62190 64766 62242 64818
rect 62638 64766 62690 64818
rect 63422 64766 63474 64818
rect 68014 64766 68066 64818
rect 72158 64766 72210 64818
rect 114830 64766 114882 64818
rect 116958 64766 117010 64818
rect 45950 64654 46002 64706
rect 46734 64654 46786 64706
rect 55358 64654 55410 64706
rect 57822 64654 57874 64706
rect 58830 64654 58882 64706
rect 60622 64654 60674 64706
rect 63646 64654 63698 64706
rect 64094 64654 64146 64706
rect 65326 64654 65378 64706
rect 65998 64654 66050 64706
rect 68462 64654 68514 64706
rect 69358 64654 69410 64706
rect 46510 64542 46562 64594
rect 47854 64542 47906 64594
rect 48190 64542 48242 64594
rect 48414 64542 48466 64594
rect 57934 64542 57986 64594
rect 58942 64542 58994 64594
rect 66446 64542 66498 64594
rect 66670 64542 66722 64594
rect 67678 64542 67730 64594
rect 69694 64542 69746 64594
rect 69918 64542 69970 64594
rect 70478 64542 70530 64594
rect 70590 64542 70642 64594
rect 70702 64542 70754 64594
rect 116174 64542 116226 64594
rect 1822 64430 1874 64482
rect 47294 64430 47346 64482
rect 47966 64430 48018 64482
rect 49198 64430 49250 64482
rect 49646 64430 49698 64482
rect 50206 64430 50258 64482
rect 50654 64430 50706 64482
rect 54238 64430 54290 64482
rect 55694 64430 55746 64482
rect 65438 64430 65490 64482
rect 66334 64430 66386 64482
rect 67118 64430 67170 64482
rect 69582 64430 69634 64482
rect 71262 64430 71314 64482
rect 71710 64430 71762 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 81278 64262 81330 64314
rect 81382 64262 81434 64314
rect 81486 64262 81538 64314
rect 111998 64262 112050 64314
rect 112102 64262 112154 64314
rect 112206 64262 112258 64314
rect 53454 64094 53506 64146
rect 54126 64094 54178 64146
rect 56702 64094 56754 64146
rect 58382 64094 58434 64146
rect 63086 64094 63138 64146
rect 65550 64094 65602 64146
rect 66558 64094 66610 64146
rect 68126 64094 68178 64146
rect 68686 64094 68738 64146
rect 70702 64094 70754 64146
rect 1934 63982 1986 64034
rect 47966 63982 48018 64034
rect 49646 63982 49698 64034
rect 62750 63982 62802 64034
rect 65662 63982 65714 64034
rect 67342 63982 67394 64034
rect 48638 63870 48690 63922
rect 50766 63870 50818 63922
rect 51214 63870 51266 63922
rect 55358 63870 55410 63922
rect 55806 63870 55858 63922
rect 57598 63870 57650 63922
rect 59054 63870 59106 63922
rect 59838 63870 59890 63922
rect 64206 63870 64258 63922
rect 64766 63870 64818 63922
rect 65326 63870 65378 63922
rect 67678 63870 67730 63922
rect 69470 63870 69522 63922
rect 70478 63870 70530 63922
rect 71150 63870 71202 63922
rect 3278 63758 3330 63810
rect 45838 63758 45890 63810
rect 49534 63758 49586 63810
rect 50430 63758 50482 63810
rect 50542 63758 50594 63810
rect 54238 63758 54290 63810
rect 54910 63758 54962 63810
rect 58494 63758 58546 63810
rect 61966 63758 62018 63810
rect 63646 63758 63698 63810
rect 63758 63758 63810 63810
rect 66222 63758 66274 63810
rect 67454 63758 67506 63810
rect 69022 63758 69074 63810
rect 49870 63646 49922 63698
rect 54350 63646 54402 63698
rect 58158 63646 58210 63698
rect 63982 63646 64034 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 96638 63478 96690 63530
rect 96742 63478 96794 63530
rect 96846 63478 96898 63530
rect 51774 63310 51826 63362
rect 51998 63310 52050 63362
rect 63198 63310 63250 63362
rect 3278 63198 3330 63250
rect 48638 63198 48690 63250
rect 51998 63198 52050 63250
rect 54238 63198 54290 63250
rect 56366 63198 56418 63250
rect 57374 63198 57426 63250
rect 57822 63198 57874 63250
rect 58270 63198 58322 63250
rect 62862 63198 62914 63250
rect 68014 63198 68066 63250
rect 70142 63198 70194 63250
rect 74510 63198 74562 63250
rect 114830 63198 114882 63250
rect 47630 63086 47682 63138
rect 51550 63086 51602 63138
rect 53566 63086 53618 63138
rect 58606 63086 58658 63138
rect 58942 63086 58994 63138
rect 59166 63086 59218 63138
rect 59614 63086 59666 63138
rect 65438 63086 65490 63138
rect 65774 63086 65826 63138
rect 71598 63086 71650 63138
rect 1934 62974 1986 63026
rect 48078 62974 48130 63026
rect 50766 62974 50818 63026
rect 58494 62974 58546 63026
rect 61406 62974 61458 63026
rect 62078 62974 62130 63026
rect 62190 62974 62242 63026
rect 62414 62974 62466 63026
rect 62750 62974 62802 63026
rect 64318 62974 64370 63026
rect 66334 62974 66386 63026
rect 69358 62974 69410 63026
rect 72382 62974 72434 63026
rect 116174 62974 116226 63026
rect 58158 62862 58210 62914
rect 61854 62862 61906 62914
rect 62974 62862 63026 62914
rect 63870 62862 63922 62914
rect 68462 62862 68514 62914
rect 69470 62862 69522 62914
rect 71038 62862 71090 62914
rect 74958 62862 75010 62914
rect 117070 62862 117122 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 81278 62694 81330 62746
rect 81382 62694 81434 62746
rect 81486 62694 81538 62746
rect 111998 62694 112050 62746
rect 112102 62694 112154 62746
rect 112206 62694 112258 62746
rect 1822 62526 1874 62578
rect 50318 62526 50370 62578
rect 54686 62526 54738 62578
rect 55246 62526 55298 62578
rect 56254 62526 56306 62578
rect 63086 62526 63138 62578
rect 63758 62526 63810 62578
rect 64654 62526 64706 62578
rect 70030 62526 70082 62578
rect 72046 62526 72098 62578
rect 45838 62414 45890 62466
rect 49534 62414 49586 62466
rect 50094 62414 50146 62466
rect 55134 62414 55186 62466
rect 56702 62414 56754 62466
rect 58494 62414 58546 62466
rect 58942 62414 58994 62466
rect 73390 62414 73442 62466
rect 74174 62414 74226 62466
rect 45502 62302 45554 62354
rect 50430 62302 50482 62354
rect 50542 62302 50594 62354
rect 51102 62302 51154 62354
rect 52894 62302 52946 62354
rect 54462 62302 54514 62354
rect 55022 62302 55074 62354
rect 58046 62302 58098 62354
rect 61854 62302 61906 62354
rect 62526 62302 62578 62354
rect 63646 62302 63698 62354
rect 63870 62302 63922 62354
rect 64094 62302 64146 62354
rect 65438 62302 65490 62354
rect 65662 62302 65714 62354
rect 66782 62302 66834 62354
rect 71710 62302 71762 62354
rect 72046 62302 72098 62354
rect 72382 62302 72434 62354
rect 73502 62302 73554 62354
rect 73726 62302 73778 62354
rect 74734 62302 74786 62354
rect 48302 62190 48354 62242
rect 53342 62190 53394 62242
rect 53790 62190 53842 62242
rect 55470 62190 55522 62242
rect 55806 62190 55858 62242
rect 57598 62190 57650 62242
rect 59726 62190 59778 62242
rect 67454 62190 67506 62242
rect 69582 62190 69634 62242
rect 70478 62190 70530 62242
rect 70926 62190 70978 62242
rect 53902 62078 53954 62130
rect 65774 62078 65826 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 96638 61910 96690 61962
rect 96742 61910 96794 61962
rect 96846 61910 96898 61962
rect 54014 61742 54066 61794
rect 55918 61742 55970 61794
rect 56478 61742 56530 61794
rect 57822 61742 57874 61794
rect 58830 61742 58882 61794
rect 3614 61630 3666 61682
rect 46286 61630 46338 61682
rect 48414 61630 48466 61682
rect 48862 61630 48914 61682
rect 49310 61630 49362 61682
rect 51214 61630 51266 61682
rect 53566 61630 53618 61682
rect 55582 61630 55634 61682
rect 55918 61630 55970 61682
rect 59278 61630 59330 61682
rect 59726 61630 59778 61682
rect 62526 61630 62578 61682
rect 68350 61630 68402 61682
rect 70814 61630 70866 61682
rect 74510 61630 74562 61682
rect 80446 61630 80498 61682
rect 114830 61630 114882 61682
rect 3054 61518 3106 61570
rect 45614 61518 45666 61570
rect 66670 61518 66722 61570
rect 67454 61518 67506 61570
rect 67902 61518 67954 61570
rect 69470 61518 69522 61570
rect 69918 61518 69970 61570
rect 71710 61518 71762 61570
rect 81118 61518 81170 61570
rect 83022 61518 83074 61570
rect 1934 61406 1986 61458
rect 54350 61406 54402 61458
rect 67566 61406 67618 61458
rect 70926 61406 70978 61458
rect 72382 61406 72434 61458
rect 116174 61406 116226 61458
rect 50878 61294 50930 61346
rect 52222 61294 52274 61346
rect 52670 61294 52722 61346
rect 54126 61294 54178 61346
rect 55022 61294 55074 61346
rect 56366 61294 56418 61346
rect 56814 61294 56866 61346
rect 57598 61294 57650 61346
rect 58046 61294 58098 61346
rect 58494 61294 58546 61346
rect 58942 61294 58994 61346
rect 67342 61294 67394 61346
rect 67678 61294 67730 61346
rect 70030 61294 70082 61346
rect 70142 61294 70194 61346
rect 74958 61294 75010 61346
rect 117070 61294 117122 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 81278 61126 81330 61178
rect 81382 61126 81434 61178
rect 81486 61126 81538 61178
rect 111998 61126 112050 61178
rect 112102 61126 112154 61178
rect 112206 61126 112258 61178
rect 45726 60958 45778 61010
rect 52670 60958 52722 61010
rect 59390 60958 59442 61010
rect 60286 60958 60338 61010
rect 61518 60958 61570 61010
rect 67678 60958 67730 61010
rect 68574 60958 68626 61010
rect 69470 60958 69522 61010
rect 71934 60958 71986 61010
rect 73614 60958 73666 61010
rect 74286 60958 74338 61010
rect 46622 60846 46674 60898
rect 56366 60846 56418 60898
rect 58382 60846 58434 60898
rect 59614 60846 59666 60898
rect 59838 60846 59890 60898
rect 61742 60846 61794 60898
rect 65662 60846 65714 60898
rect 67454 60846 67506 60898
rect 68014 60846 68066 60898
rect 70366 60846 70418 60898
rect 70926 60846 70978 60898
rect 116286 60846 116338 60898
rect 46062 60734 46114 60786
rect 46510 60734 46562 60786
rect 47742 60734 47794 60786
rect 50206 60734 50258 60786
rect 53566 60734 53618 60786
rect 54014 60734 54066 60786
rect 55134 60734 55186 60786
rect 56030 60734 56082 60786
rect 58494 60734 58546 60786
rect 59166 60734 59218 60786
rect 59502 60734 59554 60786
rect 61294 60734 61346 60786
rect 61966 60734 62018 60786
rect 62414 60734 62466 60786
rect 63534 60734 63586 60786
rect 67790 60734 67842 60786
rect 69582 60734 69634 60786
rect 69806 60734 69858 60786
rect 70254 60734 70306 60786
rect 71598 60734 71650 60786
rect 71934 60734 71986 60786
rect 72270 60734 72322 60786
rect 1822 60622 1874 60674
rect 48190 60622 48242 60674
rect 49534 60622 49586 60674
rect 50318 60622 50370 60674
rect 50990 60622 51042 60674
rect 51550 60622 51602 60674
rect 52222 60622 52274 60674
rect 53006 60622 53058 60674
rect 57710 60622 57762 60674
rect 60734 60622 60786 60674
rect 62974 60622 63026 60674
rect 63758 60622 63810 60674
rect 64430 60622 64482 60674
rect 66222 60622 66274 60674
rect 66670 60622 66722 60674
rect 68686 60622 68738 60674
rect 71038 60622 71090 60674
rect 73614 60622 73666 60674
rect 114942 60622 114994 60674
rect 116846 60622 116898 60674
rect 54014 60510 54066 60562
rect 54350 60510 54402 60562
rect 55022 60510 55074 60562
rect 55358 60510 55410 60562
rect 55470 60510 55522 60562
rect 56030 60510 56082 60562
rect 58606 60510 58658 60562
rect 65438 60510 65490 60562
rect 65774 60510 65826 60562
rect 66222 60510 66274 60562
rect 66782 60510 66834 60562
rect 73390 60510 73442 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 96638 60342 96690 60394
rect 96742 60342 96794 60394
rect 96846 60342 96898 60394
rect 51214 60174 51266 60226
rect 51886 60174 51938 60226
rect 55358 60174 55410 60226
rect 58718 60174 58770 60226
rect 59502 60174 59554 60226
rect 59950 60174 60002 60226
rect 62302 60174 62354 60226
rect 63086 60174 63138 60226
rect 68014 60174 68066 60226
rect 69918 60174 69970 60226
rect 3278 60062 3330 60114
rect 47070 60062 47122 60114
rect 47966 60062 48018 60114
rect 49198 60062 49250 60114
rect 49646 60062 49698 60114
rect 53902 60062 53954 60114
rect 56478 60062 56530 60114
rect 58494 60062 58546 60114
rect 61294 60062 61346 60114
rect 61854 60062 61906 60114
rect 62302 60062 62354 60114
rect 63534 60062 63586 60114
rect 65774 60062 65826 60114
rect 67006 60062 67058 60114
rect 67454 60062 67506 60114
rect 70478 60062 70530 60114
rect 71822 60062 71874 60114
rect 48750 59950 48802 60002
rect 49758 59950 49810 60002
rect 50206 59950 50258 60002
rect 50318 59950 50370 60002
rect 50430 59950 50482 60002
rect 51886 59950 51938 60002
rect 53566 59950 53618 60002
rect 55134 59950 55186 60002
rect 55582 59950 55634 60002
rect 55918 59950 55970 60002
rect 57038 59950 57090 60002
rect 57822 59950 57874 60002
rect 59390 59950 59442 60002
rect 59726 59950 59778 60002
rect 66558 59950 66610 60002
rect 68686 59950 68738 60002
rect 69358 59950 69410 60002
rect 71374 59950 71426 60002
rect 1934 59838 1986 59890
rect 47406 59838 47458 59890
rect 52782 59838 52834 59890
rect 54910 59838 54962 59890
rect 56702 59838 56754 59890
rect 57710 59838 57762 59890
rect 62974 59838 63026 59890
rect 63310 59838 63362 59890
rect 70030 59838 70082 59890
rect 46510 59726 46562 59778
rect 48302 59726 48354 59778
rect 49534 59726 49586 59778
rect 51326 59726 51378 59778
rect 52334 59726 52386 59778
rect 54798 59726 54850 59778
rect 57486 59726 57538 59778
rect 58494 59726 58546 59778
rect 59390 59726 59442 59778
rect 60510 59726 60562 59778
rect 62862 59726 62914 59778
rect 68126 59726 68178 59778
rect 68350 59726 68402 59778
rect 69582 59726 69634 59778
rect 69806 59726 69858 59778
rect 70926 59726 70978 59778
rect 73054 59726 73106 59778
rect 114942 59726 114994 59778
rect 115278 59726 115330 59778
rect 115838 59726 115890 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 81278 59558 81330 59610
rect 81382 59558 81434 59610
rect 81486 59558 81538 59610
rect 111998 59558 112050 59610
rect 112102 59558 112154 59610
rect 112206 59558 112258 59610
rect 55022 59390 55074 59442
rect 57822 59390 57874 59442
rect 59950 59390 60002 59442
rect 60958 59390 61010 59442
rect 62862 59390 62914 59442
rect 63646 59390 63698 59442
rect 64318 59390 64370 59442
rect 66782 59390 66834 59442
rect 67566 59390 67618 59442
rect 68910 59390 68962 59442
rect 69358 59390 69410 59442
rect 69694 59390 69746 59442
rect 69918 59390 69970 59442
rect 72046 59390 72098 59442
rect 1934 59278 1986 59330
rect 49534 59278 49586 59330
rect 49758 59278 49810 59330
rect 52894 59278 52946 59330
rect 55582 59278 55634 59330
rect 57598 59278 57650 59330
rect 58494 59278 58546 59330
rect 59054 59278 59106 59330
rect 63310 59278 63362 59330
rect 66110 59278 66162 59330
rect 48750 59166 48802 59218
rect 53566 59166 53618 59218
rect 55918 59166 55970 59218
rect 56366 59166 56418 59218
rect 57486 59166 57538 59218
rect 58718 59166 58770 59218
rect 59614 59166 59666 59218
rect 59950 59166 60002 59218
rect 60286 59166 60338 59218
rect 61182 59166 61234 59218
rect 62078 59166 62130 59218
rect 62750 59166 62802 59218
rect 63086 59166 63138 59218
rect 69470 59166 69522 59218
rect 70142 59166 70194 59218
rect 70590 59166 70642 59218
rect 3278 59054 3330 59106
rect 49646 59054 49698 59106
rect 50766 59054 50818 59106
rect 54462 59054 54514 59106
rect 58942 59054 58994 59106
rect 61630 59054 61682 59106
rect 63534 59054 63586 59106
rect 63982 59054 64034 59106
rect 65326 59054 65378 59106
rect 65886 59054 65938 59106
rect 66222 59054 66274 59106
rect 67118 59054 67170 59106
rect 68014 59054 68066 59106
rect 68462 59054 68514 59106
rect 71038 59054 71090 59106
rect 71486 59054 71538 59106
rect 54686 58942 54738 58994
rect 60846 58942 60898 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 96638 58774 96690 58826
rect 96742 58774 96794 58826
rect 96846 58774 96898 58826
rect 54574 58606 54626 58658
rect 56814 58606 56866 58658
rect 59390 58606 59442 58658
rect 59614 58606 59666 58658
rect 62190 58606 62242 58658
rect 62526 58606 62578 58658
rect 63982 58606 64034 58658
rect 64206 58606 64258 58658
rect 65326 58606 65378 58658
rect 67566 58606 67618 58658
rect 68126 58606 68178 58658
rect 68350 58606 68402 58658
rect 1822 58494 1874 58546
rect 49086 58494 49138 58546
rect 52222 58494 52274 58546
rect 52782 58494 52834 58546
rect 56030 58494 56082 58546
rect 63086 58494 63138 58546
rect 63646 58494 63698 58546
rect 67678 58494 67730 58546
rect 68126 58494 68178 58546
rect 68574 58494 68626 58546
rect 69358 58494 69410 58546
rect 70926 58494 70978 58546
rect 114830 58494 114882 58546
rect 48414 58382 48466 58434
rect 55806 58382 55858 58434
rect 56254 58382 56306 58434
rect 58046 58382 58098 58434
rect 58270 58382 58322 58434
rect 58942 58382 58994 58434
rect 59166 58382 59218 58434
rect 67230 58382 67282 58434
rect 69582 58382 69634 58434
rect 70030 58382 70082 58434
rect 70702 58382 70754 58434
rect 53454 58270 53506 58322
rect 53790 58270 53842 58322
rect 54462 58270 54514 58322
rect 55582 58270 55634 58322
rect 56030 58270 56082 58322
rect 57822 58270 57874 58322
rect 58382 58270 58434 58322
rect 63758 58270 63810 58322
rect 64878 58270 64930 58322
rect 65774 58270 65826 58322
rect 69806 58270 69858 58322
rect 116174 58270 116226 58322
rect 51326 58158 51378 58210
rect 54574 58158 54626 58210
rect 56926 58158 56978 58210
rect 57038 58158 57090 58210
rect 59054 58158 59106 58210
rect 60398 58158 60450 58210
rect 61630 58158 61682 58210
rect 62414 58158 62466 58210
rect 64542 58158 64594 58210
rect 65326 58158 65378 58210
rect 66222 58158 66274 58210
rect 70366 58158 70418 58210
rect 71038 58158 71090 58210
rect 71262 58158 71314 58210
rect 71710 58158 71762 58210
rect 117070 58158 117122 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 81278 57990 81330 58042
rect 81382 57990 81434 58042
rect 81486 57990 81538 58042
rect 111998 57990 112050 58042
rect 112102 57990 112154 58042
rect 112206 57990 112258 58042
rect 51998 57822 52050 57874
rect 52446 57822 52498 57874
rect 56030 57822 56082 57874
rect 56702 57822 56754 57874
rect 62862 57822 62914 57874
rect 70814 57822 70866 57874
rect 49534 57710 49586 57762
rect 54350 57710 54402 57762
rect 57598 57710 57650 57762
rect 60622 57710 60674 57762
rect 63982 57710 64034 57762
rect 70702 57710 70754 57762
rect 117070 57710 117122 57762
rect 49870 57598 49922 57650
rect 52894 57598 52946 57650
rect 57486 57598 57538 57650
rect 59502 57598 59554 57650
rect 62302 57598 62354 57650
rect 63646 57598 63698 57650
rect 64094 57598 64146 57650
rect 64430 57598 64482 57650
rect 64654 57598 64706 57650
rect 65774 57598 65826 57650
rect 69134 57598 69186 57650
rect 69470 57598 69522 57650
rect 69694 57598 69746 57650
rect 70254 57598 70306 57650
rect 70478 57598 70530 57650
rect 117294 57598 117346 57650
rect 47854 57486 47906 57538
rect 48414 57486 48466 57538
rect 48750 57486 48802 57538
rect 50542 57486 50594 57538
rect 50990 57486 51042 57538
rect 51438 57486 51490 57538
rect 53454 57486 53506 57538
rect 54686 57486 54738 57538
rect 55246 57486 55298 57538
rect 55582 57486 55634 57538
rect 60174 57486 60226 57538
rect 61854 57486 61906 57538
rect 63310 57486 63362 57538
rect 63534 57486 63586 57538
rect 66446 57486 66498 57538
rect 68574 57486 68626 57538
rect 69582 57486 69634 57538
rect 71150 57486 71202 57538
rect 71598 57486 71650 57538
rect 116510 57486 116562 57538
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 96638 57206 96690 57258
rect 96742 57206 96794 57258
rect 96846 57206 96898 57258
rect 41134 57038 41186 57090
rect 41470 57038 41522 57090
rect 65326 57038 65378 57090
rect 41134 56926 41186 56978
rect 56702 56926 56754 56978
rect 58046 56926 58098 56978
rect 58494 56926 58546 56978
rect 58942 56926 58994 56978
rect 59278 56926 59330 56978
rect 59838 56926 59890 56978
rect 59950 56926 60002 56978
rect 61966 56926 62018 56978
rect 62638 56926 62690 56978
rect 64430 56926 64482 56978
rect 65550 56926 65602 56978
rect 66222 56926 66274 56978
rect 67006 56926 67058 56978
rect 69246 56926 69298 56978
rect 70926 56926 70978 56978
rect 73054 56926 73106 56978
rect 3054 56814 3106 56866
rect 41694 56814 41746 56866
rect 45950 56814 46002 56866
rect 47406 56814 47458 56866
rect 48526 56814 48578 56866
rect 52670 56814 52722 56866
rect 53902 56814 53954 56866
rect 57262 56814 57314 56866
rect 57598 56814 57650 56866
rect 63982 56814 64034 56866
rect 64318 56814 64370 56866
rect 67902 56814 67954 56866
rect 70254 56814 70306 56866
rect 1934 56702 1986 56754
rect 42254 56702 42306 56754
rect 49198 56702 49250 56754
rect 54574 56702 54626 56754
rect 66670 56702 66722 56754
rect 3502 56590 3554 56642
rect 46174 56590 46226 56642
rect 46958 56590 47010 56642
rect 47966 56590 48018 56642
rect 51438 56590 51490 56642
rect 52222 56590 52274 56642
rect 57374 56590 57426 56642
rect 60062 56590 60114 56642
rect 60734 56590 60786 56642
rect 61518 56590 61570 56642
rect 65550 56590 65602 56642
rect 66894 56590 66946 56642
rect 67454 56590 67506 56642
rect 68574 56590 68626 56642
rect 73502 56590 73554 56642
rect 118078 56590 118130 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 111998 56422 112050 56474
rect 112102 56422 112154 56474
rect 112206 56422 112258 56474
rect 50094 56254 50146 56306
rect 53790 56254 53842 56306
rect 55022 56254 55074 56306
rect 57934 56254 57986 56306
rect 58606 56254 58658 56306
rect 60174 56254 60226 56306
rect 62414 56254 62466 56306
rect 64318 56254 64370 56306
rect 65438 56254 65490 56306
rect 67790 56254 67842 56306
rect 68462 56254 68514 56306
rect 68574 56254 68626 56306
rect 68686 56254 68738 56306
rect 47070 56142 47122 56194
rect 49646 56142 49698 56194
rect 51102 56142 51154 56194
rect 54462 56142 54514 56194
rect 55358 56142 55410 56194
rect 56142 56142 56194 56194
rect 59054 56142 59106 56194
rect 59726 56142 59778 56194
rect 63534 56142 63586 56194
rect 63758 56142 63810 56194
rect 80334 56142 80386 56194
rect 114494 56142 114546 56194
rect 47854 56030 47906 56082
rect 48862 56030 48914 56082
rect 50206 56030 50258 56082
rect 50542 56030 50594 56082
rect 52334 56030 52386 56082
rect 54910 56030 54962 56082
rect 55134 56030 55186 56082
rect 55918 56030 55970 56082
rect 56478 56030 56530 56082
rect 57598 56030 57650 56082
rect 59278 56030 59330 56082
rect 59502 56030 59554 56082
rect 60846 56030 60898 56082
rect 61294 56030 61346 56082
rect 66558 56030 66610 56082
rect 66670 56030 66722 56082
rect 66782 56030 66834 56082
rect 67118 56030 67170 56082
rect 68350 56030 68402 56082
rect 68910 56030 68962 56082
rect 70142 56030 70194 56082
rect 79438 56030 79490 56082
rect 79998 56030 80050 56082
rect 114942 56030 114994 56082
rect 44942 55918 44994 55970
rect 48302 55918 48354 55970
rect 49870 55918 49922 55970
rect 51438 55918 51490 55970
rect 51886 55918 51938 55970
rect 52894 55918 52946 55970
rect 53678 55918 53730 55970
rect 54686 55918 54738 55970
rect 56366 55918 56418 55970
rect 61742 55918 61794 55970
rect 62862 55918 62914 55970
rect 63646 55918 63698 55970
rect 65774 55918 65826 55970
rect 67342 55918 67394 55970
rect 67790 55918 67842 55970
rect 69582 55918 69634 55970
rect 70366 55918 70418 55970
rect 71038 55918 71090 55970
rect 71486 55918 71538 55970
rect 71934 55918 71986 55970
rect 115838 55918 115890 55970
rect 50094 55806 50146 55858
rect 50766 55806 50818 55858
rect 51886 55806 51938 55858
rect 53118 55806 53170 55858
rect 53454 55806 53506 55858
rect 53790 55806 53842 55858
rect 59166 55806 59218 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 40910 55470 40962 55522
rect 46398 55470 46450 55522
rect 49646 55470 49698 55522
rect 49982 55470 50034 55522
rect 55022 55470 55074 55522
rect 67790 55470 67842 55522
rect 68238 55470 68290 55522
rect 40014 55358 40066 55410
rect 52558 55358 52610 55410
rect 54126 55358 54178 55410
rect 56814 55358 56866 55410
rect 57486 55358 57538 55410
rect 58942 55358 58994 55410
rect 59390 55358 59442 55410
rect 60062 55358 60114 55410
rect 61294 55358 61346 55410
rect 62078 55358 62130 55410
rect 64206 55358 64258 55410
rect 64654 55358 64706 55410
rect 65550 55358 65602 55410
rect 65998 55358 66050 55410
rect 67342 55358 67394 55410
rect 67790 55358 67842 55410
rect 68574 55358 68626 55410
rect 115838 55358 115890 55410
rect 40798 55246 40850 55298
rect 46734 55246 46786 55298
rect 47518 55246 47570 55298
rect 49198 55246 49250 55298
rect 50542 55246 50594 55298
rect 51214 55246 51266 55298
rect 51550 55246 51602 55298
rect 52334 55246 52386 55298
rect 52782 55246 52834 55298
rect 53678 55246 53730 55298
rect 53902 55246 53954 55298
rect 54686 55246 54738 55298
rect 54910 55246 54962 55298
rect 55134 55246 55186 55298
rect 57934 55246 57986 55298
rect 59166 55246 59218 55298
rect 59502 55246 59554 55298
rect 61854 55246 61906 55298
rect 62302 55246 62354 55298
rect 62526 55246 62578 55298
rect 62862 55246 62914 55298
rect 68238 55246 68290 55298
rect 69694 55246 69746 55298
rect 70030 55246 70082 55298
rect 70366 55246 70418 55298
rect 70590 55246 70642 55298
rect 71486 55246 71538 55298
rect 114942 55246 114994 55298
rect 47294 55134 47346 55186
rect 50990 55134 51042 55186
rect 52110 55134 52162 55186
rect 53454 55134 53506 55186
rect 58270 55134 58322 55186
rect 62974 55134 63026 55186
rect 69582 55134 69634 55186
rect 71038 55134 71090 55186
rect 1822 55022 1874 55074
rect 39678 55022 39730 55074
rect 40686 55022 40738 55074
rect 45838 55022 45890 55074
rect 48190 55022 48242 55074
rect 48638 55022 48690 55074
rect 49758 55022 49810 55074
rect 51438 55022 51490 55074
rect 54574 55022 54626 55074
rect 55246 55022 55298 55074
rect 55918 55022 55970 55074
rect 56254 55022 56306 55074
rect 58158 55022 58210 55074
rect 59054 55022 59106 55074
rect 60622 55022 60674 55074
rect 62302 55022 62354 55074
rect 63534 55022 63586 55074
rect 65102 55022 65154 55074
rect 66446 55022 66498 55074
rect 69470 55022 69522 55074
rect 70366 55022 70418 55074
rect 71934 55022 71986 55074
rect 114382 55022 114434 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 111998 54854 112050 54906
rect 112102 54854 112154 54906
rect 112206 54854 112258 54906
rect 40798 54686 40850 54738
rect 41694 54686 41746 54738
rect 45726 54686 45778 54738
rect 46510 54686 46562 54738
rect 47854 54686 47906 54738
rect 48862 54686 48914 54738
rect 51886 54686 51938 54738
rect 53006 54686 53058 54738
rect 53902 54686 53954 54738
rect 56702 54686 56754 54738
rect 59166 54686 59218 54738
rect 64430 54686 64482 54738
rect 68686 54686 68738 54738
rect 41582 54574 41634 54626
rect 41806 54574 41858 54626
rect 46174 54574 46226 54626
rect 49534 54574 49586 54626
rect 51438 54574 51490 54626
rect 51774 54574 51826 54626
rect 63646 54574 63698 54626
rect 63870 54574 63922 54626
rect 66558 54574 66610 54626
rect 67902 54574 67954 54626
rect 68126 54574 68178 54626
rect 89966 54574 90018 54626
rect 47406 54462 47458 54514
rect 49870 54462 49922 54514
rect 50206 54462 50258 54514
rect 51214 54462 51266 54514
rect 51774 54462 51826 54514
rect 52222 54462 52274 54514
rect 54574 54462 54626 54514
rect 55022 54462 55074 54514
rect 57598 54462 57650 54514
rect 57822 54462 57874 54514
rect 58494 54462 58546 54514
rect 59390 54462 59442 54514
rect 59950 54462 60002 54514
rect 69806 54462 69858 54514
rect 89630 54462 89682 54514
rect 40350 54350 40402 54402
rect 47070 54350 47122 54402
rect 48414 54350 48466 54402
rect 49982 54350 50034 54402
rect 50878 54350 50930 54402
rect 52894 54350 52946 54402
rect 54350 54350 54402 54402
rect 55806 54350 55858 54402
rect 56254 54350 56306 54402
rect 60734 54350 60786 54402
rect 62974 54350 63026 54402
rect 65438 54350 65490 54402
rect 67342 54350 67394 54402
rect 69134 54350 69186 54402
rect 70478 54350 70530 54402
rect 72606 54350 72658 54402
rect 73278 54350 73330 54402
rect 88510 54350 88562 54402
rect 45838 54238 45890 54290
rect 46622 54238 46674 54290
rect 51998 54238 52050 54290
rect 54798 54238 54850 54290
rect 55470 54238 55522 54290
rect 56142 54238 56194 54290
rect 56926 54238 56978 54290
rect 59054 54238 59106 54290
rect 63982 54238 64034 54290
rect 68238 54238 68290 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 49646 53902 49698 53954
rect 59614 53902 59666 53954
rect 61294 53902 61346 53954
rect 61854 53902 61906 53954
rect 66894 53902 66946 53954
rect 67006 53902 67058 53954
rect 70366 53902 70418 53954
rect 46846 53790 46898 53842
rect 48750 53790 48802 53842
rect 54014 53790 54066 53842
rect 59278 53790 59330 53842
rect 63982 53790 64034 53842
rect 68126 53790 68178 53842
rect 70142 53790 70194 53842
rect 45950 53678 46002 53730
rect 48414 53678 48466 53730
rect 49422 53678 49474 53730
rect 49758 53678 49810 53730
rect 50206 53678 50258 53730
rect 50990 53678 51042 53730
rect 51886 53678 51938 53730
rect 58718 53678 58770 53730
rect 60510 53678 60562 53730
rect 61742 53678 61794 53730
rect 62638 53678 62690 53730
rect 63310 53678 63362 53730
rect 67230 53678 67282 53730
rect 67342 53678 67394 53730
rect 70030 53678 70082 53730
rect 71262 53678 71314 53730
rect 45390 53566 45442 53618
rect 48190 53566 48242 53618
rect 48638 53566 48690 53618
rect 49198 53566 49250 53618
rect 50542 53566 50594 53618
rect 51662 53566 51714 53618
rect 51774 53566 51826 53618
rect 62190 53566 62242 53618
rect 68014 53566 68066 53618
rect 46398 53454 46450 53506
rect 47294 53454 47346 53506
rect 47630 53454 47682 53506
rect 49646 53454 49698 53506
rect 52334 53454 52386 53506
rect 59502 53454 59554 53506
rect 60062 53454 60114 53506
rect 61294 53454 61346 53506
rect 66222 53454 66274 53506
rect 68238 53454 68290 53506
rect 69246 53454 69298 53506
rect 70926 53454 70978 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 111998 53286 112050 53338
rect 112102 53286 112154 53338
rect 112206 53286 112258 53338
rect 33966 53118 34018 53170
rect 42478 53118 42530 53170
rect 45726 53118 45778 53170
rect 51326 53118 51378 53170
rect 54686 53118 54738 53170
rect 55582 53118 55634 53170
rect 57934 53118 57986 53170
rect 58494 53118 58546 53170
rect 59390 53118 59442 53170
rect 61854 53118 61906 53170
rect 66222 53118 66274 53170
rect 43150 53006 43202 53058
rect 43374 53006 43426 53058
rect 51886 53006 51938 53058
rect 54014 53006 54066 53058
rect 58046 53006 58098 53058
rect 60510 53006 60562 53058
rect 68574 53006 68626 53058
rect 116286 53006 116338 53058
rect 33742 52894 33794 52946
rect 48750 52894 48802 52946
rect 49758 52894 49810 52946
rect 50430 52894 50482 52946
rect 53678 52894 53730 52946
rect 56030 52894 56082 52946
rect 56254 52894 56306 52946
rect 56702 52894 56754 52946
rect 58158 52894 58210 52946
rect 58718 52894 58770 52946
rect 61406 52894 61458 52946
rect 63870 52894 63922 52946
rect 65774 52894 65826 52946
rect 66334 52894 66386 52946
rect 66446 52894 66498 52946
rect 67790 52894 67842 52946
rect 34414 52782 34466 52834
rect 42030 52782 42082 52834
rect 43262 52782 43314 52834
rect 47966 52782 48018 52834
rect 52334 52782 52386 52834
rect 52782 52782 52834 52834
rect 53230 52782 53282 52834
rect 54798 52782 54850 52834
rect 57374 52782 57426 52834
rect 57710 52782 57762 52834
rect 59278 52782 59330 52834
rect 60062 52782 60114 52834
rect 60958 52782 61010 52834
rect 62302 52782 62354 52834
rect 63310 52782 63362 52834
rect 64542 52782 64594 52834
rect 65326 52782 65378 52834
rect 65550 52782 65602 52834
rect 65774 52782 65826 52834
rect 66894 52782 66946 52834
rect 70702 52782 70754 52834
rect 114942 52782 114994 52834
rect 116846 52782 116898 52834
rect 49870 52670 49922 52722
rect 52334 52670 52386 52722
rect 53342 52670 53394 52722
rect 54910 52670 54962 52722
rect 56478 52670 56530 52722
rect 59614 52670 59666 52722
rect 60734 52670 60786 52722
rect 61406 52670 61458 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 46622 52334 46674 52386
rect 48190 52334 48242 52386
rect 48638 52334 48690 52386
rect 49198 52334 49250 52386
rect 49534 52334 49586 52386
rect 50094 52334 50146 52386
rect 50430 52334 50482 52386
rect 52222 52334 52274 52386
rect 55918 52334 55970 52386
rect 56366 52334 56418 52386
rect 60286 52334 60338 52386
rect 60622 52334 60674 52386
rect 62414 52334 62466 52386
rect 67790 52334 67842 52386
rect 3278 52222 3330 52274
rect 46062 52222 46114 52274
rect 47294 52222 47346 52274
rect 47742 52222 47794 52274
rect 48190 52222 48242 52274
rect 51998 52222 52050 52274
rect 56814 52222 56866 52274
rect 57262 52222 57314 52274
rect 57710 52222 57762 52274
rect 58158 52222 58210 52274
rect 63086 52222 63138 52274
rect 64430 52222 64482 52274
rect 65102 52222 65154 52274
rect 67230 52222 67282 52274
rect 68574 52222 68626 52274
rect 69694 52222 69746 52274
rect 73502 52222 73554 52274
rect 74062 52222 74114 52274
rect 46398 52110 46450 52162
rect 48638 52110 48690 52162
rect 51102 52110 51154 52162
rect 54462 52110 54514 52162
rect 54798 52110 54850 52162
rect 55470 52110 55522 52162
rect 55694 52110 55746 52162
rect 61406 52110 61458 52162
rect 63982 52110 64034 52162
rect 65214 52110 65266 52162
rect 66670 52110 66722 52162
rect 67006 52110 67058 52162
rect 69246 52110 69298 52162
rect 70702 52110 70754 52162
rect 1934 51998 1986 52050
rect 54238 51998 54290 52050
rect 59390 51998 59442 52050
rect 64990 51998 65042 52050
rect 65438 51998 65490 52050
rect 71374 51998 71426 52050
rect 46958 51886 47010 51938
rect 49310 51886 49362 51938
rect 50318 51886 50370 51938
rect 50990 51886 51042 51938
rect 52558 51886 52610 51938
rect 53790 51886 53842 51938
rect 58830 51886 58882 51938
rect 58942 51886 58994 51938
rect 59054 51886 59106 51938
rect 59166 51886 59218 51938
rect 60510 51886 60562 51938
rect 67902 51886 67954 51938
rect 68014 51886 68066 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 111998 51718 112050 51770
rect 112102 51718 112154 51770
rect 112206 51718 112258 51770
rect 1822 51550 1874 51602
rect 48414 51550 48466 51602
rect 49646 51550 49698 51602
rect 51550 51550 51602 51602
rect 56366 51550 56418 51602
rect 58046 51550 58098 51602
rect 58830 51550 58882 51602
rect 59390 51550 59442 51602
rect 66222 51550 66274 51602
rect 66782 51550 66834 51602
rect 67230 51550 67282 51602
rect 67566 51550 67618 51602
rect 71150 51550 71202 51602
rect 73278 51550 73330 51602
rect 45054 51438 45106 51490
rect 47518 51438 47570 51490
rect 47742 51438 47794 51490
rect 52894 51438 52946 51490
rect 53902 51438 53954 51490
rect 56254 51438 56306 51490
rect 56478 51438 56530 51490
rect 57486 51438 57538 51490
rect 58606 51438 58658 51490
rect 64542 51438 64594 51490
rect 65438 51438 65490 51490
rect 69470 51438 69522 51490
rect 70926 51438 70978 51490
rect 72046 51438 72098 51490
rect 50878 51326 50930 51378
rect 53118 51326 53170 51378
rect 54014 51326 54066 51378
rect 57710 51326 57762 51378
rect 58942 51326 58994 51378
rect 60286 51326 60338 51378
rect 64094 51326 64146 51378
rect 65774 51326 65826 51378
rect 68126 51326 68178 51378
rect 68910 51326 68962 51378
rect 71150 51326 71202 51378
rect 71486 51326 71538 51378
rect 72158 51326 72210 51378
rect 72382 51326 72434 51378
rect 45502 51214 45554 51266
rect 46062 51214 46114 51266
rect 46510 51214 46562 51266
rect 46958 51214 47010 51266
rect 47630 51214 47682 51266
rect 48302 51214 48354 51266
rect 49982 51214 50034 51266
rect 61070 51214 61122 51266
rect 63310 51214 63362 51266
rect 69918 51214 69970 51266
rect 70478 51214 70530 51266
rect 73726 51214 73778 51266
rect 45614 51102 45666 51154
rect 46510 51102 46562 51154
rect 50542 51102 50594 51154
rect 50878 51102 50930 51154
rect 51438 51102 51490 51154
rect 51774 51102 51826 51154
rect 52446 51102 52498 51154
rect 68798 51102 68850 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 53342 50766 53394 50818
rect 53566 50766 53618 50818
rect 54238 50766 54290 50818
rect 61518 50766 61570 50818
rect 67342 50766 67394 50818
rect 68798 50766 68850 50818
rect 45502 50654 45554 50706
rect 49198 50654 49250 50706
rect 50430 50654 50482 50706
rect 52670 50654 52722 50706
rect 53566 50654 53618 50706
rect 55470 50654 55522 50706
rect 56478 50654 56530 50706
rect 58494 50654 58546 50706
rect 59390 50654 59442 50706
rect 60510 50654 60562 50706
rect 64430 50654 64482 50706
rect 65214 50654 65266 50706
rect 67230 50654 67282 50706
rect 68238 50654 68290 50706
rect 68574 50654 68626 50706
rect 72270 50654 72322 50706
rect 115502 50654 115554 50706
rect 48302 50542 48354 50594
rect 50654 50542 50706 50594
rect 50878 50542 50930 50594
rect 51214 50542 51266 50594
rect 52222 50542 52274 50594
rect 54910 50542 54962 50594
rect 56142 50542 56194 50594
rect 58606 50542 58658 50594
rect 59726 50542 59778 50594
rect 59950 50542 60002 50594
rect 62190 50542 62242 50594
rect 63758 50542 63810 50594
rect 64542 50542 64594 50594
rect 65662 50542 65714 50594
rect 66558 50542 66610 50594
rect 67790 50542 67842 50594
rect 69358 50542 69410 50594
rect 72718 50542 72770 50594
rect 116174 50542 116226 50594
rect 117294 50542 117346 50594
rect 47630 50430 47682 50482
rect 50206 50430 50258 50482
rect 51662 50430 51714 50482
rect 51886 50430 51938 50482
rect 54350 50430 54402 50482
rect 55246 50430 55298 50482
rect 61630 50430 61682 50482
rect 64318 50430 64370 50482
rect 70142 50430 70194 50482
rect 117070 50430 117122 50482
rect 49758 50318 49810 50370
rect 50766 50318 50818 50370
rect 51550 50318 51602 50370
rect 54238 50318 54290 50370
rect 63422 50318 63474 50370
rect 64766 50318 64818 50370
rect 66670 50318 66722 50370
rect 66894 50318 66946 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 111998 50150 112050 50202
rect 112102 50150 112154 50202
rect 112206 50150 112258 50202
rect 45838 49982 45890 50034
rect 46398 49982 46450 50034
rect 47070 49982 47122 50034
rect 47966 49982 48018 50034
rect 48750 49982 48802 50034
rect 50430 49982 50482 50034
rect 53230 49982 53282 50034
rect 54574 49982 54626 50034
rect 63198 49982 63250 50034
rect 64430 49982 64482 50034
rect 70030 49982 70082 50034
rect 116846 49982 116898 50034
rect 47406 49870 47458 49922
rect 50878 49870 50930 49922
rect 52110 49870 52162 49922
rect 52334 49870 52386 49922
rect 53678 49870 53730 49922
rect 54350 49870 54402 49922
rect 55022 49870 55074 49922
rect 60622 49870 60674 49922
rect 64206 49870 64258 49922
rect 72046 49870 72098 49922
rect 72270 49870 72322 49922
rect 45502 49758 45554 49810
rect 46734 49758 46786 49810
rect 47070 49758 47122 49810
rect 50206 49758 50258 49810
rect 50430 49758 50482 49810
rect 50542 49758 50594 49810
rect 54238 49758 54290 49810
rect 56366 49758 56418 49810
rect 56814 49758 56866 49810
rect 57822 49758 57874 49810
rect 63982 49758 64034 49810
rect 66782 49758 66834 49810
rect 68126 49758 68178 49810
rect 69806 49758 69858 49810
rect 70030 49758 70082 49810
rect 70366 49758 70418 49810
rect 70926 49758 70978 49810
rect 45054 49646 45106 49698
rect 48414 49646 48466 49698
rect 49534 49646 49586 49698
rect 51550 49646 51602 49698
rect 52110 49646 52162 49698
rect 52782 49646 52834 49698
rect 64094 49646 64146 49698
rect 65326 49646 65378 49698
rect 65774 49646 65826 49698
rect 66894 49646 66946 49698
rect 68574 49646 68626 49698
rect 69022 49646 69074 49698
rect 71486 49646 71538 49698
rect 72270 49646 72322 49698
rect 73278 49646 73330 49698
rect 67230 49534 67282 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 51102 49198 51154 49250
rect 70590 49198 70642 49250
rect 70926 49198 70978 49250
rect 46510 49086 46562 49138
rect 46958 49086 47010 49138
rect 47854 49086 47906 49138
rect 48414 49086 48466 49138
rect 48862 49086 48914 49138
rect 50318 49086 50370 49138
rect 52670 49086 52722 49138
rect 53454 49086 53506 49138
rect 54126 49086 54178 49138
rect 58830 49086 58882 49138
rect 61518 49086 61570 49138
rect 62974 49086 63026 49138
rect 64654 49086 64706 49138
rect 68014 49086 68066 49138
rect 68350 49086 68402 49138
rect 69582 49086 69634 49138
rect 70590 49086 70642 49138
rect 71822 49086 71874 49138
rect 115502 49086 115554 49138
rect 49310 48974 49362 49026
rect 49534 48974 49586 49026
rect 49646 48974 49698 49026
rect 49982 48974 50034 49026
rect 50542 48974 50594 49026
rect 53902 48974 53954 49026
rect 55246 48974 55298 49026
rect 56478 48974 56530 49026
rect 57486 48974 57538 49026
rect 57710 48974 57762 49026
rect 59950 48974 60002 49026
rect 61630 48974 61682 49026
rect 62078 48974 62130 49026
rect 62862 48974 62914 49026
rect 63198 48974 63250 49026
rect 63870 48974 63922 49026
rect 116174 48974 116226 49026
rect 46062 48862 46114 48914
rect 52110 48862 52162 48914
rect 54238 48862 54290 48914
rect 55134 48862 55186 48914
rect 55358 48862 55410 48914
rect 60062 48862 60114 48914
rect 61406 48862 61458 48914
rect 63086 48862 63138 48914
rect 1822 48750 1874 48802
rect 45726 48750 45778 48802
rect 47406 48750 47458 48802
rect 50318 48750 50370 48802
rect 51214 48750 51266 48802
rect 51326 48750 51378 48802
rect 51998 48750 52050 48802
rect 55806 48750 55858 48802
rect 56926 48750 56978 48802
rect 58046 48750 58098 48802
rect 62750 48750 62802 48802
rect 66894 48750 66946 48802
rect 67454 48750 67506 48802
rect 71038 48750 71090 48802
rect 116958 48750 117010 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 111998 48582 112050 48634
rect 112102 48582 112154 48634
rect 112206 48582 112258 48634
rect 45278 48414 45330 48466
rect 48862 48414 48914 48466
rect 56702 48414 56754 48466
rect 58718 48414 58770 48466
rect 64206 48414 64258 48466
rect 65886 48414 65938 48466
rect 67118 48414 67170 48466
rect 67678 48414 67730 48466
rect 117070 48414 117122 48466
rect 46734 48302 46786 48354
rect 47070 48302 47122 48354
rect 47966 48302 48018 48354
rect 49646 48302 49698 48354
rect 49870 48302 49922 48354
rect 51550 48302 51602 48354
rect 53006 48302 53058 48354
rect 58158 48302 58210 48354
rect 58830 48302 58882 48354
rect 61742 48302 61794 48354
rect 67230 48302 67282 48354
rect 68462 48302 68514 48354
rect 47294 48190 47346 48242
rect 49534 48190 49586 48242
rect 52110 48190 52162 48242
rect 52446 48190 52498 48242
rect 55246 48190 55298 48242
rect 57598 48190 57650 48242
rect 59166 48190 59218 48242
rect 59614 48190 59666 48242
rect 60510 48190 60562 48242
rect 61294 48190 61346 48242
rect 61518 48190 61570 48242
rect 63086 48190 63138 48242
rect 63310 48190 63362 48242
rect 63982 48190 64034 48242
rect 64318 48190 64370 48242
rect 66110 48190 66162 48242
rect 67342 48190 67394 48242
rect 67902 48190 67954 48242
rect 68798 48190 68850 48242
rect 70142 48190 70194 48242
rect 116174 48190 116226 48242
rect 117294 48190 117346 48242
rect 45726 48078 45778 48130
rect 46286 48078 46338 48130
rect 46846 48078 46898 48130
rect 47854 48078 47906 48130
rect 50766 48078 50818 48130
rect 54798 48078 54850 48130
rect 55694 48078 55746 48130
rect 56142 48078 56194 48130
rect 58382 48078 58434 48130
rect 60398 48078 60450 48130
rect 61406 48078 61458 48130
rect 66670 48078 66722 48130
rect 67006 48078 67058 48130
rect 68686 48078 68738 48130
rect 69246 48078 69298 48130
rect 69694 48078 69746 48130
rect 70590 48078 70642 48130
rect 115502 48078 115554 48130
rect 48190 47966 48242 48018
rect 58606 47966 58658 48018
rect 63198 47966 63250 48018
rect 65774 47966 65826 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 54014 47630 54066 47682
rect 55022 47630 55074 47682
rect 55358 47630 55410 47682
rect 56030 47630 56082 47682
rect 57374 47630 57426 47682
rect 57710 47630 57762 47682
rect 58270 47630 58322 47682
rect 59614 47630 59666 47682
rect 62190 47630 62242 47682
rect 62974 47630 63026 47682
rect 3278 47518 3330 47570
rect 45502 47518 45554 47570
rect 47630 47518 47682 47570
rect 48974 47518 49026 47570
rect 51102 47518 51154 47570
rect 52670 47518 52722 47570
rect 53790 47518 53842 47570
rect 54574 47518 54626 47570
rect 56254 47518 56306 47570
rect 57710 47518 57762 47570
rect 59950 47518 60002 47570
rect 60398 47518 60450 47570
rect 63086 47518 63138 47570
rect 67678 47518 67730 47570
rect 68350 47518 68402 47570
rect 71150 47518 71202 47570
rect 73278 47518 73330 47570
rect 73726 47518 73778 47570
rect 2606 47406 2658 47458
rect 48414 47406 48466 47458
rect 51774 47406 51826 47458
rect 55582 47406 55634 47458
rect 55918 47406 55970 47458
rect 57374 47406 57426 47458
rect 59054 47406 59106 47458
rect 61294 47406 61346 47458
rect 61630 47406 61682 47458
rect 62302 47406 62354 47458
rect 63310 47406 63362 47458
rect 67006 47406 67058 47458
rect 70366 47406 70418 47458
rect 117294 47406 117346 47458
rect 56478 47294 56530 47346
rect 58718 47294 58770 47346
rect 58830 47294 58882 47346
rect 66222 47294 66274 47346
rect 67566 47294 67618 47346
rect 69246 47294 69298 47346
rect 117070 47294 117122 47346
rect 2830 47182 2882 47234
rect 53790 47182 53842 47234
rect 55022 47182 55074 47234
rect 56030 47182 56082 47234
rect 59838 47182 59890 47234
rect 61518 47182 61570 47234
rect 63982 47182 64034 47234
rect 67790 47182 67842 47234
rect 69806 47182 69858 47234
rect 116286 47182 116338 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 111998 47014 112050 47066
rect 112102 47014 112154 47066
rect 112206 47014 112258 47066
rect 46846 46846 46898 46898
rect 47518 46846 47570 46898
rect 48750 46846 48802 46898
rect 54350 46846 54402 46898
rect 56590 46846 56642 46898
rect 57374 46846 57426 46898
rect 58270 46846 58322 46898
rect 64094 46846 64146 46898
rect 65326 46846 65378 46898
rect 65774 46846 65826 46898
rect 66670 46846 66722 46898
rect 47294 46734 47346 46786
rect 55806 46734 55858 46786
rect 56030 46734 56082 46786
rect 59950 46734 60002 46786
rect 62638 46734 62690 46786
rect 63198 46734 63250 46786
rect 66222 46734 66274 46786
rect 68686 46734 68738 46786
rect 118078 46734 118130 46786
rect 2830 46622 2882 46674
rect 47630 46622 47682 46674
rect 47854 46622 47906 46674
rect 49870 46622 49922 46674
rect 50542 46622 50594 46674
rect 59278 46622 59330 46674
rect 62862 46622 62914 46674
rect 62974 46622 63026 46674
rect 63086 46622 63138 46674
rect 63758 46622 63810 46674
rect 64094 46622 64146 46674
rect 64318 46622 64370 46674
rect 68014 46622 68066 46674
rect 1934 46510 1986 46562
rect 48414 46510 48466 46562
rect 49982 46510 50034 46562
rect 51326 46510 51378 46562
rect 53454 46510 53506 46562
rect 54686 46510 54738 46562
rect 55134 46510 55186 46562
rect 58606 46510 58658 46562
rect 62078 46510 62130 46562
rect 67230 46510 67282 46562
rect 70814 46510 70866 46562
rect 55694 46398 55746 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 50654 46062 50706 46114
rect 52446 46062 52498 46114
rect 52670 46062 52722 46114
rect 59614 46062 59666 46114
rect 59838 46062 59890 46114
rect 45614 45950 45666 46002
rect 47742 45950 47794 46002
rect 50206 45950 50258 46002
rect 50878 45950 50930 46002
rect 52222 45950 52274 46002
rect 52670 45950 52722 46002
rect 53678 45950 53730 46002
rect 55358 45950 55410 46002
rect 60622 45950 60674 46002
rect 67230 45950 67282 46002
rect 115502 45950 115554 46002
rect 3054 45838 3106 45890
rect 48526 45838 48578 45890
rect 54126 45838 54178 45890
rect 54574 45838 54626 45890
rect 58606 45838 58658 45890
rect 58942 45838 58994 45890
rect 61406 45838 61458 45890
rect 116174 45838 116226 45890
rect 1934 45726 1986 45778
rect 63870 45726 63922 45778
rect 68014 45726 68066 45778
rect 3502 45614 3554 45666
rect 49198 45614 49250 45666
rect 49646 45614 49698 45666
rect 50878 45614 50930 45666
rect 51550 45614 51602 45666
rect 57598 45614 57650 45666
rect 58718 45614 58770 45666
rect 59614 45614 59666 45666
rect 60174 45614 60226 45666
rect 67566 45614 67618 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 42926 45278 42978 45330
rect 47742 45278 47794 45330
rect 48638 45278 48690 45330
rect 49422 45278 49474 45330
rect 50990 45278 51042 45330
rect 51438 45278 51490 45330
rect 52446 45278 52498 45330
rect 54910 45278 54962 45330
rect 56366 45278 56418 45330
rect 56814 45278 56866 45330
rect 57486 45278 57538 45330
rect 61630 45278 61682 45330
rect 61966 45278 62018 45330
rect 64206 45278 64258 45330
rect 64542 45278 64594 45330
rect 116510 45278 116562 45330
rect 117070 45278 117122 45330
rect 42142 45166 42194 45218
rect 42478 45166 42530 45218
rect 51998 45166 52050 45218
rect 53678 45166 53730 45218
rect 58830 45166 58882 45218
rect 59502 45166 59554 45218
rect 65774 45166 65826 45218
rect 117406 45166 117458 45218
rect 46958 45054 47010 45106
rect 47518 45054 47570 45106
rect 58270 45054 58322 45106
rect 58494 45054 58546 45106
rect 59278 45054 59330 45106
rect 59614 45054 59666 45106
rect 63422 45054 63474 45106
rect 50542 44942 50594 44994
rect 53230 44942 53282 44994
rect 54126 44942 54178 44994
rect 54462 44942 54514 44994
rect 55358 44942 55410 44994
rect 55918 44942 55970 44994
rect 58382 44942 58434 44994
rect 60062 44942 60114 44994
rect 60510 44942 60562 44994
rect 60958 44942 61010 44994
rect 62750 44942 62802 44994
rect 65326 44942 65378 44994
rect 66446 44942 66498 44994
rect 66894 44942 66946 44994
rect 47854 44830 47906 44882
rect 54238 44830 54290 44882
rect 55022 44830 55074 44882
rect 60622 44830 60674 44882
rect 60958 44830 61010 44882
rect 62078 44830 62130 44882
rect 62974 44830 63026 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 49086 44494 49138 44546
rect 50318 44494 50370 44546
rect 52110 44494 52162 44546
rect 61966 44494 62018 44546
rect 49086 44382 49138 44434
rect 50430 44382 50482 44434
rect 54238 44382 54290 44434
rect 55918 44382 55970 44434
rect 56702 44382 56754 44434
rect 57374 44382 57426 44434
rect 59502 44382 59554 44434
rect 65102 44382 65154 44434
rect 67902 44382 67954 44434
rect 49982 44270 50034 44322
rect 51886 44270 51938 44322
rect 55022 44270 55074 44322
rect 60286 44270 60338 44322
rect 61294 44270 61346 44322
rect 62414 44270 62466 44322
rect 65662 44270 65714 44322
rect 66110 44270 66162 44322
rect 66894 44270 66946 44322
rect 67230 44270 67282 44322
rect 51326 44158 51378 44210
rect 53678 44158 53730 44210
rect 53790 44158 53842 44210
rect 53902 44158 53954 44210
rect 54798 44158 54850 44210
rect 55358 44158 55410 44210
rect 62974 44158 63026 44210
rect 64206 44158 64258 44210
rect 67454 44158 67506 44210
rect 48078 44046 48130 44098
rect 49534 44046 49586 44098
rect 50878 44046 50930 44098
rect 52446 44046 52498 44098
rect 53454 44046 53506 44098
rect 55134 44046 55186 44098
rect 61630 44046 61682 44098
rect 61854 44046 61906 44098
rect 67006 44046 67058 44098
rect 67118 44046 67170 44098
rect 68462 44046 68514 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 59950 43710 60002 43762
rect 61630 43710 61682 43762
rect 64542 43710 64594 43762
rect 68238 43710 68290 43762
rect 52894 43598 52946 43650
rect 54238 43598 54290 43650
rect 57486 43598 57538 43650
rect 63086 43598 63138 43650
rect 63534 43598 63586 43650
rect 66222 43598 66274 43650
rect 116286 43598 116338 43650
rect 50430 43486 50482 43538
rect 50766 43486 50818 43538
rect 51886 43486 51938 43538
rect 53566 43486 53618 43538
rect 58494 43486 58546 43538
rect 58942 43486 58994 43538
rect 60286 43486 60338 43538
rect 61966 43486 62018 43538
rect 62302 43486 62354 43538
rect 62414 43486 62466 43538
rect 62750 43486 62802 43538
rect 65326 43486 65378 43538
rect 87278 43486 87330 43538
rect 48302 43374 48354 43426
rect 48862 43374 48914 43426
rect 49870 43374 49922 43426
rect 51998 43374 52050 43426
rect 52446 43374 52498 43426
rect 56366 43374 56418 43426
rect 58046 43374 58098 43426
rect 63982 43374 64034 43426
rect 82350 43374 82402 43426
rect 87838 43374 87890 43426
rect 114942 43374 114994 43426
rect 116846 43374 116898 43426
rect 59950 43262 60002 43314
rect 60062 43262 60114 43314
rect 60510 43262 60562 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 48750 42814 48802 42866
rect 50430 42814 50482 42866
rect 50878 42814 50930 42866
rect 52222 42814 52274 42866
rect 54910 42814 54962 42866
rect 55358 42814 55410 42866
rect 55918 42814 55970 42866
rect 56366 42814 56418 42866
rect 56702 42814 56754 42866
rect 57262 42814 57314 42866
rect 58830 42814 58882 42866
rect 60622 42814 60674 42866
rect 61742 42814 61794 42866
rect 62190 42814 62242 42866
rect 62750 42814 62802 42866
rect 63198 42814 63250 42866
rect 64430 42814 64482 42866
rect 48190 42702 48242 42754
rect 49534 42702 49586 42754
rect 49870 42702 49922 42754
rect 50206 42702 50258 42754
rect 51550 42702 51602 42754
rect 51774 42702 51826 42754
rect 52110 42702 52162 42754
rect 52558 42702 52610 42754
rect 57934 42702 57986 42754
rect 58270 42702 58322 42754
rect 59166 42702 59218 42754
rect 59614 42702 59666 42754
rect 59950 42702 60002 42754
rect 48974 42590 49026 42642
rect 49758 42590 49810 42642
rect 53454 42590 53506 42642
rect 53678 42590 53730 42642
rect 54238 42590 54290 42642
rect 57710 42590 57762 42642
rect 59502 42590 59554 42642
rect 61406 42590 61458 42642
rect 61630 42590 61682 42642
rect 63534 42590 63586 42642
rect 63982 42590 64034 42642
rect 47742 42478 47794 42530
rect 50542 42478 50594 42530
rect 51438 42478 51490 42530
rect 52670 42478 52722 42530
rect 53566 42478 53618 42530
rect 58046 42478 58098 42530
rect 58158 42478 58210 42530
rect 59390 42478 59442 42530
rect 60062 42478 60114 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 56814 42142 56866 42194
rect 63982 42142 64034 42194
rect 58158 42030 58210 42082
rect 61742 42030 61794 42082
rect 54798 41918 54850 41970
rect 55246 41918 55298 41970
rect 55694 41918 55746 41970
rect 57934 41918 57986 41970
rect 59390 41918 59442 41970
rect 60958 41918 61010 41970
rect 114382 41918 114434 41970
rect 114942 41918 114994 41970
rect 48302 41806 48354 41858
rect 48750 41806 48802 41858
rect 52782 41806 52834 41858
rect 57374 41806 57426 41858
rect 59278 41806 59330 41858
rect 60398 41806 60450 41858
rect 115838 41806 115890 41858
rect 58270 41694 58322 41746
rect 59502 41694 59554 41746
rect 60062 41694 60114 41746
rect 60398 41694 60450 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 57150 41358 57202 41410
rect 57710 41358 57762 41410
rect 3278 41246 3330 41298
rect 49198 41246 49250 41298
rect 52670 41246 52722 41298
rect 54238 41246 54290 41298
rect 56366 41246 56418 41298
rect 57150 41246 57202 41298
rect 58718 41246 58770 41298
rect 59502 41246 59554 41298
rect 61406 41246 61458 41298
rect 61518 41246 61570 41298
rect 115502 41246 115554 41298
rect 47518 41134 47570 41186
rect 49870 41134 49922 41186
rect 53454 41134 53506 41186
rect 59054 41134 59106 41186
rect 116174 41134 116226 41186
rect 1934 41022 1986 41074
rect 50542 41022 50594 41074
rect 47742 40910 47794 40962
rect 57598 40910 57650 40962
rect 58158 40910 58210 40962
rect 60174 40910 60226 40962
rect 60622 40910 60674 40962
rect 61630 40910 61682 40962
rect 62190 40910 62242 40962
rect 62750 40910 62802 40962
rect 116958 40910 117010 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 49422 40574 49474 40626
rect 50878 40574 50930 40626
rect 51550 40574 51602 40626
rect 52334 40574 52386 40626
rect 53118 40574 53170 40626
rect 54126 40574 54178 40626
rect 54462 40574 54514 40626
rect 61966 40574 62018 40626
rect 117070 40574 117122 40626
rect 1710 40462 1762 40514
rect 47966 40462 48018 40514
rect 53678 40462 53730 40514
rect 61182 40462 61234 40514
rect 116286 40462 116338 40514
rect 48750 40350 48802 40402
rect 52670 40350 52722 40402
rect 61518 40350 61570 40402
rect 62414 40350 62466 40402
rect 117294 40350 117346 40402
rect 45838 40238 45890 40290
rect 50654 40238 50706 40290
rect 50990 40238 51042 40290
rect 61294 40238 61346 40290
rect 115166 40238 115218 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 48078 39790 48130 39842
rect 3614 39678 3666 39730
rect 47406 39678 47458 39730
rect 48414 39678 48466 39730
rect 49870 39678 49922 39730
rect 51326 39678 51378 39730
rect 53342 39678 53394 39730
rect 117070 39678 117122 39730
rect 3054 39566 3106 39618
rect 49198 39566 49250 39618
rect 1934 39454 1986 39506
rect 48974 39454 49026 39506
rect 50206 39454 50258 39506
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 61070 39006 61122 39058
rect 63422 39006 63474 39058
rect 53790 38894 53842 38946
rect 62862 38894 62914 38946
rect 63870 38894 63922 38946
rect 118078 38894 118130 38946
rect 53566 38782 53618 38834
rect 62078 38782 62130 38834
rect 62638 38782 62690 38834
rect 61742 38558 61794 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 52782 38110 52834 38162
rect 54238 38110 54290 38162
rect 56366 38110 56418 38162
rect 64318 38110 64370 38162
rect 3054 37998 3106 38050
rect 53454 37998 53506 38050
rect 61406 37998 61458 38050
rect 1934 37886 1986 37938
rect 62190 37886 62242 37938
rect 3502 37774 3554 37826
rect 60622 37774 60674 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 54238 37438 54290 37490
rect 56030 37438 56082 37490
rect 61854 37438 61906 37490
rect 1934 37326 1986 37378
rect 54910 37326 54962 37378
rect 55134 37326 55186 37378
rect 54574 37214 54626 37266
rect 61630 37214 61682 37266
rect 3278 37102 3330 37154
rect 53566 37102 53618 37154
rect 56366 37102 56418 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 3278 36542 3330 36594
rect 114830 36542 114882 36594
rect 2158 36318 2210 36370
rect 116174 36318 116226 36370
rect 117070 36206 117122 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 1822 35870 1874 35922
rect 2158 35758 2210 35810
rect 114494 35646 114546 35698
rect 114942 35646 114994 35698
rect 115838 35534 115890 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 3278 34974 3330 35026
rect 45838 34862 45890 34914
rect 116174 34862 116226 34914
rect 1934 34750 1986 34802
rect 58270 34750 58322 34802
rect 46062 34638 46114 34690
rect 57710 34638 57762 34690
rect 58606 34638 58658 34690
rect 115950 34638 116002 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 47182 34190 47234 34242
rect 115950 34190 116002 34242
rect 3054 34078 3106 34130
rect 47966 34078 48018 34130
rect 115166 34078 115218 34130
rect 1934 33966 1986 34018
rect 3614 33966 3666 34018
rect 45054 33966 45106 34018
rect 48414 33966 48466 34018
rect 114606 33966 114658 34018
rect 118078 33966 118130 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 46062 33518 46114 33570
rect 1822 33406 1874 33458
rect 45390 33406 45442 33458
rect 46398 33406 46450 33458
rect 47742 33406 47794 33458
rect 115502 33406 115554 33458
rect 48190 33294 48242 33346
rect 116062 33294 116114 33346
rect 46622 33182 46674 33234
rect 46958 33182 47010 33234
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 116062 32734 116114 32786
rect 1934 32622 1986 32674
rect 114942 32622 114994 32674
rect 116622 32622 116674 32674
rect 117182 32622 117234 32674
rect 3278 32398 3330 32450
rect 115390 32398 115442 32450
rect 116398 32286 116450 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 1822 31838 1874 31890
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 116174 30942 116226 30994
rect 115502 30830 115554 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 116174 30382 116226 30434
rect 116510 30382 116562 30434
rect 3278 30270 3330 30322
rect 69358 30158 69410 30210
rect 114382 30158 114434 30210
rect 114942 30158 114994 30210
rect 115502 30158 115554 30210
rect 1934 30046 1986 30098
rect 72270 30046 72322 30098
rect 117070 30046 117122 30098
rect 117406 30046 117458 30098
rect 75070 29934 75122 29986
rect 116286 29934 116338 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 1822 29598 1874 29650
rect 49422 29598 49474 29650
rect 47742 29374 47794 29426
rect 48526 29150 48578 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 45502 28478 45554 28530
rect 45838 28366 45890 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 48190 28030 48242 28082
rect 46958 27918 47010 27970
rect 47742 27806 47794 27858
rect 44830 27694 44882 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 45726 27246 45778 27298
rect 46062 27246 46114 27298
rect 3278 27134 3330 27186
rect 47406 27134 47458 27186
rect 47854 27134 47906 27186
rect 115502 27134 115554 27186
rect 46846 27022 46898 27074
rect 116174 27022 116226 27074
rect 1934 26910 1986 26962
rect 44718 26910 44770 26962
rect 46622 26910 46674 26962
rect 117070 26910 117122 26962
rect 117406 26910 117458 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 63198 26462 63250 26514
rect 116734 26462 116786 26514
rect 1710 26350 1762 26402
rect 58830 26350 58882 26402
rect 62750 26238 62802 26290
rect 114382 26238 114434 26290
rect 114942 26238 114994 26290
rect 2158 26126 2210 26178
rect 115838 26126 115890 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 3278 25566 3330 25618
rect 45614 25454 45666 25506
rect 1934 25342 1986 25394
rect 45838 25230 45890 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 48078 24894 48130 24946
rect 46846 24782 46898 24834
rect 3054 24670 3106 24722
rect 47630 24670 47682 24722
rect 1934 24558 1986 24610
rect 3502 24558 3554 24610
rect 44718 24558 44770 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 45726 24110 45778 24162
rect 77870 24110 77922 24162
rect 78430 24110 78482 24162
rect 77870 23998 77922 24050
rect 46062 23886 46114 23938
rect 46846 23886 46898 23938
rect 44718 23774 44770 23826
rect 46622 23774 46674 23826
rect 47406 23774 47458 23826
rect 47854 23662 47906 23714
rect 78318 23662 78370 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 116622 23326 116674 23378
rect 45838 23214 45890 23266
rect 77870 23214 77922 23266
rect 79102 23214 79154 23266
rect 79662 23214 79714 23266
rect 117070 23214 117122 23266
rect 3054 23102 3106 23154
rect 45614 23102 45666 23154
rect 77646 23102 77698 23154
rect 78542 23102 78594 23154
rect 78878 23102 78930 23154
rect 117294 23102 117346 23154
rect 1934 22990 1986 23042
rect 3502 22990 3554 23042
rect 80222 22990 80274 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 48190 22430 48242 22482
rect 76526 22430 76578 22482
rect 78318 22430 78370 22482
rect 80446 22430 80498 22482
rect 115502 22430 115554 22482
rect 46398 22318 46450 22370
rect 47182 22318 47234 22370
rect 77534 22318 77586 22370
rect 116174 22318 116226 22370
rect 1934 22206 1986 22258
rect 46958 22206 47010 22258
rect 47742 22206 47794 22258
rect 91758 22206 91810 22258
rect 4398 22094 4450 22146
rect 45502 22094 45554 22146
rect 46062 22094 46114 22146
rect 92094 22094 92146 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 48414 21758 48466 21810
rect 44494 21646 44546 21698
rect 47182 21646 47234 21698
rect 91982 21646 92034 21698
rect 3054 21534 3106 21586
rect 44270 21534 44322 21586
rect 47966 21534 48018 21586
rect 91310 21534 91362 21586
rect 1934 21422 1986 21474
rect 3614 21422 3666 21474
rect 45054 21422 45106 21474
rect 90638 21422 90690 21474
rect 94110 21422 94162 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 91198 20974 91250 21026
rect 1822 20862 1874 20914
rect 40238 20862 40290 20914
rect 45502 20862 45554 20914
rect 47630 20862 47682 20914
rect 48974 20862 49026 20914
rect 93102 20862 93154 20914
rect 39790 20750 39842 20802
rect 48302 20750 48354 20802
rect 91534 20750 91586 20802
rect 92206 20750 92258 20802
rect 39454 20638 39506 20690
rect 92318 20638 92370 20690
rect 90078 20526 90130 20578
rect 90526 20526 90578 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 45502 20078 45554 20130
rect 46062 20078 46114 20130
rect 46958 20078 47010 20130
rect 47182 19966 47234 20018
rect 48302 19966 48354 20018
rect 47742 19854 47794 19906
rect 46398 19742 46450 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 115502 19294 115554 19346
rect 116174 19182 116226 19234
rect 117406 19182 117458 19234
rect 117070 19070 117122 19122
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 116734 18622 116786 18674
rect 1822 18510 1874 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 1822 17390 1874 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 118078 16942 118130 16994
rect 3054 16830 3106 16882
rect 3502 16830 3554 16882
rect 1934 16718 1986 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 54462 15374 54514 15426
rect 114494 15374 114546 15426
rect 54126 15262 54178 15314
rect 114942 15262 114994 15314
rect 53678 15150 53730 15202
rect 115838 15150 115890 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 115838 14590 115890 14642
rect 114494 14478 114546 14530
rect 114942 14478 114994 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 116286 12238 116338 12290
rect 2830 12126 2882 12178
rect 1934 12014 1986 12066
rect 114942 12014 114994 12066
rect 116846 12014 116898 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 3278 11454 3330 11506
rect 2606 11342 2658 11394
rect 2830 11230 2882 11282
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 3054 10558 3106 10610
rect 1934 10446 1986 10498
rect 3502 10446 3554 10498
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 115502 9886 115554 9938
rect 116174 9774 116226 9826
rect 117294 9774 117346 9826
rect 117070 9662 117122 9714
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 116734 9214 116786 9266
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 63870 8318 63922 8370
rect 115838 8318 115890 8370
rect 64430 8206 64482 8258
rect 114494 8206 114546 8258
rect 114942 8206 114994 8258
rect 64766 7982 64818 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 1822 7534 1874 7586
rect 116174 7422 116226 7474
rect 2382 7310 2434 7362
rect 115502 7310 115554 7362
rect 116734 7310 116786 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 114830 6750 114882 6802
rect 3054 6638 3106 6690
rect 1934 6526 1986 6578
rect 116174 6526 116226 6578
rect 117070 6526 117122 6578
rect 117406 6526 117458 6578
rect 3614 6414 3666 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 112366 6078 112418 6130
rect 116286 5966 116338 6018
rect 3054 5854 3106 5906
rect 3502 5854 3554 5906
rect 113150 5854 113202 5906
rect 1934 5742 1986 5794
rect 5182 5742 5234 5794
rect 42030 5742 42082 5794
rect 48078 5742 48130 5794
rect 113822 5742 113874 5794
rect 114942 5742 114994 5794
rect 116846 5742 116898 5794
rect 117294 5742 117346 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 5630 5182 5682 5234
rect 6078 5182 6130 5234
rect 43262 5182 43314 5234
rect 46174 5182 46226 5234
rect 47294 5182 47346 5234
rect 49198 5182 49250 5234
rect 50318 5182 50370 5234
rect 112814 5182 112866 5234
rect 114830 5182 114882 5234
rect 2830 5070 2882 5122
rect 4846 5070 4898 5122
rect 25230 5070 25282 5122
rect 26350 5070 26402 5122
rect 26910 5070 26962 5122
rect 41582 5070 41634 5122
rect 46622 5070 46674 5122
rect 59838 5070 59890 5122
rect 63982 5070 64034 5122
rect 1934 4958 1986 5010
rect 3726 4958 3778 5010
rect 40686 4958 40738 5010
rect 42366 4958 42418 5010
rect 48414 4958 48466 5010
rect 54798 4958 54850 5010
rect 55246 4958 55298 5010
rect 99150 4958 99202 5010
rect 111358 4958 111410 5010
rect 111918 4958 111970 5010
rect 114158 4958 114210 5010
rect 116174 4958 116226 5010
rect 42702 4846 42754 4898
rect 43710 4846 43762 4898
rect 48750 4846 48802 4898
rect 54462 4846 54514 4898
rect 99486 4846 99538 4898
rect 99934 4846 99986 4898
rect 101390 4846 101442 4898
rect 112254 4846 112306 4898
rect 117070 4846 117122 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 6526 4510 6578 4562
rect 9662 4510 9714 4562
rect 10558 4510 10610 4562
rect 11902 4510 11954 4562
rect 15374 4510 15426 4562
rect 28142 4510 28194 4562
rect 32846 4510 32898 4562
rect 46846 4510 46898 4562
rect 49422 4510 49474 4562
rect 57374 4510 57426 4562
rect 62974 4510 63026 4562
rect 65326 4510 65378 4562
rect 68686 4510 68738 4562
rect 76526 4510 76578 4562
rect 78318 4510 78370 4562
rect 80558 4510 80610 4562
rect 81678 4510 81730 4562
rect 104302 4510 104354 4562
rect 1934 4398 1986 4450
rect 5630 4398 5682 4450
rect 5966 4398 6018 4450
rect 11454 4398 11506 4450
rect 18510 4398 18562 4450
rect 44046 4398 44098 4450
rect 45950 4398 46002 4450
rect 46286 4398 46338 4450
rect 49982 4398 50034 4450
rect 50654 4398 50706 4450
rect 50990 4398 51042 4450
rect 53454 4398 53506 4450
rect 61070 4398 61122 4450
rect 67790 4398 67842 4450
rect 68126 4398 68178 4450
rect 71822 4398 71874 4450
rect 76974 4398 77026 4450
rect 77310 4398 77362 4450
rect 87950 4398 88002 4450
rect 93998 4398 94050 4450
rect 99374 4398 99426 4450
rect 101166 4398 101218 4450
rect 103518 4398 103570 4450
rect 103854 4398 103906 4450
rect 116286 4398 116338 4450
rect 117070 4398 117122 4450
rect 117406 4398 117458 4450
rect 4958 4286 5010 4338
rect 8206 4286 8258 4338
rect 11230 4286 11282 4338
rect 14926 4286 14978 4338
rect 27694 4286 27746 4338
rect 32174 4286 32226 4338
rect 43150 4286 43202 4338
rect 48526 4286 48578 4338
rect 51550 4286 51602 4338
rect 56590 4286 56642 4338
rect 59502 4286 59554 4338
rect 63422 4286 63474 4338
rect 73390 4286 73442 4338
rect 78878 4286 78930 4338
rect 83470 4286 83522 4338
rect 95006 4286 95058 4338
rect 100942 4286 100994 4338
rect 101726 4286 101778 4338
rect 112366 4286 112418 4338
rect 113150 4286 113202 4338
rect 3278 4174 3330 4226
rect 3950 4174 4002 4226
rect 7086 4174 7138 4226
rect 8766 4174 8818 4226
rect 13806 4174 13858 4226
rect 17950 4174 18002 4226
rect 19630 4174 19682 4226
rect 21198 4174 21250 4226
rect 21534 4174 21586 4226
rect 26574 4174 26626 4226
rect 31278 4174 31330 4226
rect 36542 4174 36594 4226
rect 37662 4174 37714 4226
rect 42254 4174 42306 4226
rect 45390 4174 45442 4226
rect 47406 4174 47458 4226
rect 52222 4174 52274 4226
rect 54686 4174 54738 4226
rect 55470 4174 55522 4226
rect 58382 4174 58434 4226
rect 60062 4174 60114 4226
rect 64094 4174 64146 4226
rect 70366 4174 70418 4226
rect 70814 4174 70866 4226
rect 74062 4174 74114 4226
rect 75742 4174 75794 4226
rect 79550 4174 79602 4226
rect 82350 4174 82402 4226
rect 86494 4174 86546 4226
rect 86942 4174 86994 4226
rect 92542 4174 92594 4226
rect 92990 4174 93042 4226
rect 95678 4174 95730 4226
rect 97918 4174 97970 4226
rect 98366 4174 98418 4226
rect 100270 4174 100322 4226
rect 102398 4174 102450 4226
rect 111694 4174 111746 4226
rect 113822 4174 113874 4226
rect 114942 4174 114994 4226
rect 117854 4174 117906 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 4958 3614 5010 3666
rect 6414 3614 6466 3666
rect 7982 3614 8034 3666
rect 12238 3614 12290 3666
rect 16494 3614 16546 3666
rect 20638 3614 20690 3666
rect 22654 3614 22706 3666
rect 26798 3614 26850 3666
rect 31054 3614 31106 3666
rect 35534 3614 35586 3666
rect 39118 3614 39170 3666
rect 43262 3614 43314 3666
rect 46510 3614 46562 3666
rect 49534 3614 49586 3666
rect 54686 3614 54738 3666
rect 59502 3614 59554 3666
rect 63758 3614 63810 3666
rect 65438 3614 65490 3666
rect 69470 3614 69522 3666
rect 73166 3614 73218 3666
rect 74174 3614 74226 3666
rect 78206 3614 78258 3666
rect 81678 3614 81730 3666
rect 84142 3614 84194 3666
rect 88510 3614 88562 3666
rect 91982 3614 92034 3666
rect 94782 3614 94834 3666
rect 96350 3614 96402 3666
rect 100494 3614 100546 3666
rect 104414 3614 104466 3666
rect 111582 3614 111634 3666
rect 115502 3614 115554 3666
rect 117406 3614 117458 3666
rect 2830 3502 2882 3554
rect 5966 3502 6018 3554
rect 8766 3502 8818 3554
rect 10670 3502 10722 3554
rect 11566 3502 11618 3554
rect 36318 3502 36370 3554
rect 48862 3502 48914 3554
rect 51662 3502 51714 3554
rect 64990 3502 65042 3554
rect 77534 3502 77586 3554
rect 80894 3502 80946 3554
rect 89966 3502 90018 3554
rect 99822 3502 99874 3554
rect 102622 3502 102674 3554
rect 103854 3502 103906 3554
rect 2046 3390 2098 3442
rect 3838 3390 3890 3442
rect 9774 3390 9826 3442
rect 14590 3390 14642 3442
rect 15150 3390 15202 3442
rect 19630 3390 19682 3442
rect 21534 3390 21586 3442
rect 24670 3390 24722 3442
rect 25454 3390 25506 3442
rect 29374 3390 29426 3442
rect 29934 3390 29986 3442
rect 37998 3390 38050 3442
rect 41470 3390 41522 3442
rect 42030 3390 42082 3442
rect 44270 3390 44322 3442
rect 45390 3390 45442 3442
rect 50766 3390 50818 3442
rect 53118 3390 53170 3442
rect 55806 3390 55858 3442
rect 56590 3390 56642 3442
rect 57598 3390 57650 3442
rect 58158 3390 58210 3442
rect 62750 3390 62802 3442
rect 69022 3390 69074 3442
rect 70478 3390 70530 3442
rect 75070 3390 75122 3442
rect 83470 3390 83522 3442
rect 85150 3390 85202 3442
rect 89070 3390 89122 3442
rect 91310 3390 91362 3442
rect 92990 3390 93042 3442
rect 95902 3390 95954 3442
rect 97358 3390 97410 3442
rect 101726 3390 101778 3442
rect 110910 3390 110962 3442
rect 112590 3390 112642 3442
rect 114158 3390 114210 3442
rect 114494 3390 114546 3442
rect 116510 3390 116562 3442
rect 2494 3278 2546 3330
rect 27694 3278 27746 3330
rect 28478 3278 28530 3330
rect 33182 3278 33234 3330
rect 37214 3278 37266 3330
rect 76302 3278 76354 3330
rect 80222 3278 80274 3330
rect 105534 3278 105586 3330
rect 109118 3278 109170 3330
rect 109790 3278 109842 3330
rect 118078 3278 118130 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 104302 1710 104354 1762
rect 105534 1710 105586 1762
<< metal2 >>
rect -56 119336 168 119800
rect 1288 119336 1512 119800
rect -56 119200 196 119336
rect 1288 119200 1540 119336
rect 1960 119200 2184 119800
rect 3304 119336 3528 119800
rect 3304 119200 3556 119336
rect 4648 119200 4872 119800
rect 5992 119336 6216 119800
rect 5964 119200 6216 119336
rect 6664 119200 6888 119800
rect 8008 119200 8232 119800
rect 9352 119200 9576 119800
rect 10024 119200 10248 119800
rect 11368 119336 11592 119800
rect 11368 119200 11620 119336
rect 12712 119200 12936 119800
rect 14056 119200 14280 119800
rect 14728 119200 14952 119800
rect 16072 119336 16296 119800
rect 16044 119200 16296 119336
rect 17416 119200 17640 119800
rect 18760 119336 18984 119800
rect 18760 119200 19012 119336
rect 19432 119200 19656 119800
rect 20776 119200 21000 119800
rect 22120 119336 22344 119800
rect 22092 119200 22344 119336
rect 22792 119200 23016 119800
rect 24136 119336 24360 119800
rect 24136 119200 24388 119336
rect 25480 119200 25704 119800
rect 26824 119200 27048 119800
rect 27496 119200 27720 119800
rect 28840 119336 29064 119800
rect 28812 119200 29064 119336
rect 30184 119200 30408 119800
rect 31528 119336 31752 119800
rect 32200 119336 32424 119800
rect 31500 119200 31752 119336
rect 32172 119200 32424 119336
rect 33544 119336 33768 119800
rect 34888 119336 35112 119800
rect 35560 119336 35784 119800
rect 33544 119200 33796 119336
rect 34888 119200 35140 119336
rect 140 117908 196 119200
rect 140 117842 196 117852
rect 1484 117124 1540 119200
rect 2044 118916 2100 118926
rect 1820 117908 1876 117918
rect 1708 117124 1764 117134
rect 1484 117122 1764 117124
rect 1484 117070 1710 117122
rect 1762 117070 1764 117122
rect 1484 117068 1764 117070
rect 1708 117058 1764 117068
rect 1820 115780 1876 117852
rect 1932 117122 1988 117134
rect 1932 117070 1934 117122
rect 1986 117070 1988 117122
rect 1932 116338 1988 117070
rect 1932 116286 1934 116338
rect 1986 116286 1988 116338
rect 1932 116004 1988 116286
rect 1932 115938 1988 115948
rect 1932 115780 1988 115790
rect 1820 115778 1988 115780
rect 1820 115726 1934 115778
rect 1986 115726 1988 115778
rect 1820 115724 1988 115726
rect 1932 115714 1988 115724
rect 2044 114994 2100 118860
rect 3388 116676 3444 116686
rect 3276 116564 3332 116574
rect 3388 116564 3444 116620
rect 3276 116562 3444 116564
rect 3276 116510 3278 116562
rect 3330 116510 3444 116562
rect 3276 116508 3444 116510
rect 3276 116498 3332 116508
rect 3052 116228 3108 116238
rect 3052 115666 3108 116172
rect 3500 115780 3556 119200
rect 4476 116844 4740 116854
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4476 116778 4740 116788
rect 5852 116564 5908 116574
rect 5964 116564 6020 119200
rect 5852 116562 6468 116564
rect 5852 116510 5854 116562
rect 5906 116510 6468 116562
rect 5852 116508 6468 116510
rect 5852 116498 5908 116508
rect 4060 116450 4116 116462
rect 4060 116398 4062 116450
rect 4114 116398 4116 116450
rect 3836 116228 3892 116238
rect 3836 116134 3892 116172
rect 3724 115780 3780 115790
rect 4060 115780 4116 116398
rect 6412 116338 6468 116508
rect 6412 116286 6414 116338
rect 6466 116286 6468 116338
rect 6412 116274 6468 116286
rect 7532 116562 7588 116574
rect 7532 116510 7534 116562
rect 7586 116510 7588 116562
rect 3500 115778 3780 115780
rect 3500 115726 3726 115778
rect 3778 115726 3780 115778
rect 3500 115724 3780 115726
rect 3724 115714 3780 115724
rect 3836 115724 4116 115780
rect 4732 116226 4788 116238
rect 4732 116174 4734 116226
rect 4786 116174 4788 116226
rect 4732 115780 4788 116174
rect 5740 115892 5796 115902
rect 5740 115798 5796 115836
rect 3052 115614 3054 115666
rect 3106 115614 3108 115666
rect 3052 115602 3108 115614
rect 2044 114942 2046 114994
rect 2098 114942 2100 114994
rect 2044 114930 2100 114942
rect 3164 114996 3220 115006
rect 3052 114884 3108 114894
rect 3052 114790 3108 114828
rect 2380 114660 2436 114670
rect 1932 114212 1988 114222
rect 1820 114210 1988 114212
rect 1820 114158 1934 114210
rect 1986 114158 1988 114210
rect 1820 114156 1988 114158
rect 1820 113540 1876 114156
rect 1932 114146 1988 114156
rect 1820 113426 1876 113484
rect 1820 113374 1822 113426
rect 1874 113374 1876 113426
rect 1820 113362 1876 113374
rect 1932 112420 1988 112430
rect 1932 112326 1988 112364
rect 1932 111636 1988 111646
rect 1708 111634 1988 111636
rect 1708 111582 1934 111634
rect 1986 111582 1988 111634
rect 1708 111580 1988 111582
rect 1708 111076 1764 111580
rect 1932 111570 1988 111580
rect 1708 110982 1764 111020
rect 1820 109954 1876 109966
rect 1820 109902 1822 109954
rect 1874 109902 1876 109954
rect 1820 109732 1876 109902
rect 1820 109666 1876 109676
rect 1820 107938 1876 107950
rect 1820 107886 1822 107938
rect 1874 107886 1876 107938
rect 1820 107716 1876 107886
rect 1820 107650 1876 107660
rect 1932 104578 1988 104590
rect 1932 104526 1934 104578
rect 1986 104526 1988 104578
rect 1932 104356 1988 104526
rect 1932 104290 1988 104300
rect 1932 103012 1988 103022
rect 1932 102918 1988 102956
rect 2380 102508 2436 114604
rect 2828 113204 2884 113214
rect 2828 113202 2996 113204
rect 2828 113150 2830 113202
rect 2882 113150 2996 113202
rect 2828 113148 2996 113150
rect 2828 113138 2884 113148
rect 2492 113090 2548 113102
rect 2492 113038 2494 113090
rect 2546 113038 2548 113090
rect 2492 112532 2548 113038
rect 2940 113092 2996 113148
rect 3164 113092 3220 114940
rect 3612 114996 3668 115006
rect 3612 114882 3668 114940
rect 3836 114996 3892 115724
rect 4732 115714 4788 115724
rect 4620 115668 4676 115678
rect 3836 114930 3892 114940
rect 3948 115666 4676 115668
rect 3948 115614 4622 115666
rect 4674 115614 4676 115666
rect 3948 115612 4676 115614
rect 3612 114830 3614 114882
rect 3666 114830 3668 114882
rect 3612 114818 3668 114830
rect 3724 114884 3780 114894
rect 3724 114098 3780 114828
rect 3948 114770 4004 115612
rect 4620 115602 4676 115612
rect 5292 115556 5348 115566
rect 4476 115276 4740 115286
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4476 115210 4740 115220
rect 4396 114996 4452 115006
rect 4396 114902 4452 114940
rect 5292 114996 5348 115500
rect 5292 114930 5348 114940
rect 3948 114718 3950 114770
rect 4002 114718 4004 114770
rect 3948 114706 4004 114718
rect 3724 114046 3726 114098
rect 3778 114046 3780 114098
rect 3276 113988 3332 113998
rect 3724 113988 3780 114046
rect 3276 113986 3444 113988
rect 3276 113934 3278 113986
rect 3330 113934 3444 113986
rect 3276 113932 3444 113934
rect 3276 113922 3332 113932
rect 3388 113876 3444 113932
rect 3724 113922 3780 113932
rect 3388 113810 3444 113820
rect 4476 113708 4740 113718
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4476 113642 4740 113652
rect 3276 113092 3332 113102
rect 2940 113090 3332 113092
rect 2940 113038 3278 113090
rect 3330 113038 3332 113090
rect 2940 113036 3332 113038
rect 2828 112532 2884 112542
rect 2492 112530 2884 112532
rect 2492 112478 2830 112530
rect 2882 112478 2884 112530
rect 2492 112476 2884 112478
rect 2828 112466 2884 112476
rect 2380 102452 2548 102508
rect 2268 102228 2324 102238
rect 2268 102226 2436 102228
rect 2268 102174 2270 102226
rect 2322 102174 2436 102226
rect 2268 102172 2436 102174
rect 2268 102162 2324 102172
rect 1820 101666 1876 101678
rect 1820 101614 1822 101666
rect 1874 101614 1876 101666
rect 1820 100996 1876 101614
rect 2380 101668 2436 102172
rect 2380 101574 2436 101612
rect 1820 100930 1876 100940
rect 1932 100100 1988 100110
rect 1820 100098 1988 100100
rect 1820 100046 1934 100098
rect 1986 100046 1988 100098
rect 1820 100044 1988 100046
rect 1820 99428 1876 100044
rect 1932 100034 1988 100044
rect 1820 99314 1876 99372
rect 1820 99262 1822 99314
rect 1874 99262 1876 99314
rect 1820 99250 1876 99262
rect 2492 99204 2548 102452
rect 2604 99204 2660 99214
rect 2492 99148 2604 99204
rect 2604 99110 2660 99148
rect 2828 98978 2884 98990
rect 2828 98926 2830 98978
rect 2882 98926 2884 98978
rect 2828 98418 2884 98926
rect 2828 98366 2830 98418
rect 2882 98366 2884 98418
rect 2828 98354 2884 98366
rect 1932 98308 1988 98318
rect 1932 98214 1988 98252
rect 1932 97524 1988 97534
rect 1708 97522 1988 97524
rect 1708 97470 1934 97522
rect 1986 97470 1988 97522
rect 1708 97468 1988 97470
rect 1708 96964 1764 97468
rect 1932 97458 1988 97468
rect 1708 96870 1764 96908
rect 2828 95282 2884 95294
rect 2828 95230 2830 95282
rect 2882 95230 2884 95282
rect 1932 95170 1988 95182
rect 1932 95118 1934 95170
rect 1986 95118 1988 95170
rect 1932 94948 1988 95118
rect 1932 94882 1988 94892
rect 2828 94724 2884 95230
rect 2716 94668 2884 94724
rect 2940 94724 2996 113036
rect 3276 113026 3332 113036
rect 4476 112140 4740 112150
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4476 112074 4740 112084
rect 3276 111860 3332 111870
rect 3276 111766 3332 111804
rect 4476 110572 4740 110582
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4476 110506 4740 110516
rect 4476 109004 4740 109014
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4476 108938 4740 108948
rect 4476 107436 4740 107446
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4476 107370 4740 107380
rect 4476 105868 4740 105878
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4476 105802 4740 105812
rect 3052 104690 3108 104702
rect 3052 104638 3054 104690
rect 3106 104638 3108 104690
rect 3052 104580 3108 104638
rect 3052 104514 3108 104524
rect 3612 104580 3668 104590
rect 3612 104486 3668 104524
rect 4476 104300 4740 104310
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4476 104234 4740 104244
rect 3052 103122 3108 103134
rect 3052 103070 3054 103122
rect 3106 103070 3108 103122
rect 3052 103012 3108 103070
rect 3052 102946 3108 102956
rect 3612 103012 3668 103022
rect 3612 102918 3668 102956
rect 4476 102732 4740 102742
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4476 102666 4740 102676
rect 3164 102452 3220 102462
rect 3164 102358 3220 102396
rect 4476 101164 4740 101174
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4476 101098 4740 101108
rect 3276 99876 3332 99886
rect 3276 99782 3332 99820
rect 4476 99596 4740 99606
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4476 99530 4740 99540
rect 3164 99204 3220 99214
rect 3164 98980 3220 99148
rect 3276 98980 3332 98990
rect 3164 98978 3332 98980
rect 3164 98926 3278 98978
rect 3330 98926 3332 98978
rect 3164 98924 3332 98926
rect 3164 94948 3220 98924
rect 3276 98914 3332 98924
rect 4476 98028 4740 98038
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4476 97962 4740 97972
rect 3276 97748 3332 97758
rect 3276 97654 3332 97692
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 3164 94892 3444 94948
rect 2940 94668 3332 94724
rect 2492 94388 2548 94398
rect 2716 94388 2772 94668
rect 2492 94386 2772 94388
rect 2492 94334 2494 94386
rect 2546 94334 2772 94386
rect 2492 94332 2772 94334
rect 2828 94500 2884 94510
rect 2940 94500 2996 94668
rect 3276 94610 3332 94668
rect 3276 94558 3278 94610
rect 3330 94558 3332 94610
rect 3276 94546 3332 94558
rect 2828 94498 2996 94500
rect 2828 94446 2830 94498
rect 2882 94446 2996 94498
rect 2828 94444 2996 94446
rect 2492 94322 2548 94332
rect 1932 93604 1988 93614
rect 1932 93510 1988 93548
rect 1932 92820 1988 92830
rect 1820 92372 1876 92382
rect 1932 92372 1988 92764
rect 1820 92370 1988 92372
rect 1820 92318 1822 92370
rect 1874 92318 1988 92370
rect 1820 92316 1988 92318
rect 1820 92306 1876 92316
rect 2828 90748 2884 94444
rect 3388 94388 3444 94892
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 3276 94332 3444 94388
rect 3276 94276 3332 94332
rect 3164 94220 3332 94276
rect 3052 93714 3108 93726
rect 3052 93662 3054 93714
rect 3106 93662 3108 93714
rect 3052 93604 3108 93662
rect 3052 93538 3108 93548
rect 2828 90692 2996 90748
rect 2828 90580 2884 90590
rect 2492 90578 2884 90580
rect 2492 90526 2830 90578
rect 2882 90526 2884 90578
rect 2492 90524 2884 90526
rect 1932 90466 1988 90478
rect 1932 90414 1934 90466
rect 1986 90414 1988 90466
rect 1932 90244 1988 90414
rect 1932 90178 1988 90188
rect 2492 89682 2548 90524
rect 2828 90514 2884 90524
rect 2940 90020 2996 90692
rect 3052 90020 3108 90030
rect 2940 90018 3108 90020
rect 2940 89966 3054 90018
rect 3106 89966 3108 90018
rect 2940 89964 3108 89966
rect 2828 89796 2884 89806
rect 2940 89796 2996 89964
rect 3052 89954 3108 89964
rect 2828 89794 2996 89796
rect 2828 89742 2830 89794
rect 2882 89742 2996 89794
rect 2828 89740 2996 89742
rect 2828 89730 2884 89740
rect 2492 89630 2494 89682
rect 2546 89630 2548 89682
rect 2492 89618 2548 89630
rect 1932 88900 1988 88910
rect 1932 88806 1988 88844
rect 1932 88116 1988 88126
rect 1820 87668 1876 87678
rect 1932 87668 1988 88060
rect 1820 87666 1988 87668
rect 1820 87614 1822 87666
rect 1874 87614 1988 87666
rect 1820 87612 1988 87614
rect 1820 87602 1876 87612
rect 1820 85986 1876 85998
rect 1820 85934 1822 85986
rect 1874 85934 1876 85986
rect 1820 85540 1876 85934
rect 1820 85474 1876 85484
rect 1820 84418 1876 84430
rect 1820 84366 1822 84418
rect 1874 84366 1876 84418
rect 1820 84196 1876 84366
rect 1820 84130 1876 84140
rect 2828 82740 2884 82750
rect 2492 82738 2884 82740
rect 2492 82686 2830 82738
rect 2882 82686 2884 82738
rect 2492 82684 2884 82686
rect 1932 82626 1988 82638
rect 1932 82574 1934 82626
rect 1986 82574 1988 82626
rect 1932 82180 1988 82574
rect 1932 82114 1988 82124
rect 2492 81842 2548 82684
rect 2828 82674 2884 82684
rect 2940 82180 2996 89740
rect 3052 89012 3108 89022
rect 3052 88918 3108 88956
rect 3052 82180 3108 82190
rect 2940 82178 3108 82180
rect 2940 82126 3054 82178
rect 3106 82126 3108 82178
rect 2940 82124 3108 82126
rect 2828 81956 2884 81966
rect 2940 81956 2996 82124
rect 3052 82114 3108 82124
rect 2828 81954 2996 81956
rect 2828 81902 2830 81954
rect 2882 81902 2996 81954
rect 2828 81900 2996 81902
rect 2828 81890 2884 81900
rect 2492 81790 2494 81842
rect 2546 81790 2548 81842
rect 2492 81778 2548 81790
rect 2828 80388 2884 80398
rect 2492 80386 2884 80388
rect 2492 80334 2830 80386
rect 2882 80334 2884 80386
rect 2492 80332 2884 80334
rect 1932 80274 1988 80286
rect 1932 80222 1934 80274
rect 1986 80222 1988 80274
rect 1932 80164 1988 80222
rect 1932 80098 1988 80108
rect 2492 79826 2548 80332
rect 2828 80322 2884 80332
rect 2492 79774 2494 79826
rect 2546 79774 2548 79826
rect 2492 79762 2548 79774
rect 2828 79602 2884 79614
rect 2828 79550 2830 79602
rect 2882 79550 2884 79602
rect 2828 79380 2884 79550
rect 3052 79380 3108 79390
rect 2828 79378 3108 79380
rect 2828 79326 3054 79378
rect 3106 79326 3108 79378
rect 2828 79324 3108 79326
rect 3052 79314 3108 79324
rect 3164 78988 3220 94220
rect 3612 93604 3668 93614
rect 3612 93510 3668 93548
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 3276 93044 3332 93054
rect 3276 92950 3332 92988
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 3276 90018 3332 90030
rect 3276 89966 3278 90018
rect 3330 89966 3332 90018
rect 3276 89906 3332 89966
rect 3276 89854 3278 89906
rect 3330 89854 3332 89906
rect 3276 89842 3332 89854
rect 5068 89684 5124 89694
rect 3500 89012 3556 89022
rect 3500 88918 3556 88956
rect 5068 89012 5124 89628
rect 5068 88946 5124 88956
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 3276 88340 3332 88350
rect 3276 88246 3332 88284
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 2940 78932 3220 78988
rect 3276 82178 3332 82190
rect 3276 82126 3278 82178
rect 3330 82126 3332 82178
rect 3276 82066 3332 82126
rect 3276 82014 3278 82066
rect 3330 82014 3332 82066
rect 3276 79826 3332 82014
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 3276 79774 3278 79826
rect 3330 79774 3332 79826
rect 3276 79378 3332 79774
rect 3276 79326 3278 79378
rect 3330 79326 3332 79378
rect 1932 78708 1988 78718
rect 1932 78614 1988 78652
rect 1820 77028 1876 77038
rect 1820 77026 1988 77028
rect 1820 76974 1822 77026
rect 1874 76974 1988 77026
rect 1820 76972 1988 76974
rect 1820 76962 1876 76972
rect 1932 76578 1988 76972
rect 1932 76526 1934 76578
rect 1986 76526 1988 76578
rect 1932 76132 1988 76526
rect 1932 76066 1988 76076
rect 2828 75684 2884 75694
rect 2492 75682 2884 75684
rect 2492 75630 2830 75682
rect 2882 75630 2884 75682
rect 2492 75628 2884 75630
rect 1932 75570 1988 75582
rect 1932 75518 1934 75570
rect 1986 75518 1988 75570
rect 1932 75460 1988 75518
rect 1932 75394 1988 75404
rect 2492 75122 2548 75628
rect 2828 75618 2884 75628
rect 2492 75070 2494 75122
rect 2546 75070 2548 75122
rect 2492 75058 2548 75070
rect 2828 75012 2884 75022
rect 1932 71876 1988 71886
rect 1820 71874 1988 71876
rect 1820 71822 1934 71874
rect 1986 71822 1988 71874
rect 1820 71820 1988 71822
rect 1820 71204 1876 71820
rect 1932 71810 1988 71820
rect 1820 71090 1876 71148
rect 1820 71038 1822 71090
rect 1874 71038 1876 71090
rect 1820 71026 1876 71038
rect 2828 70420 2884 74956
rect 2492 70306 2548 70318
rect 2492 70254 2494 70306
rect 2546 70254 2548 70306
rect 2492 69412 2548 70254
rect 2828 70306 2884 70364
rect 2828 70254 2830 70306
rect 2882 70254 2884 70306
rect 2828 70242 2884 70254
rect 2828 69412 2884 69422
rect 2492 69410 2884 69412
rect 2492 69358 2830 69410
rect 2882 69358 2884 69410
rect 2492 69356 2884 69358
rect 2828 69346 2884 69356
rect 1932 69300 1988 69310
rect 1932 69206 1988 69244
rect 1932 68514 1988 68526
rect 1932 68462 1934 68514
rect 1986 68462 1988 68514
rect 1932 68068 1988 68462
rect 1932 68002 1988 68012
rect 2940 67228 2996 78932
rect 3052 78818 3108 78830
rect 3052 78766 3054 78818
rect 3106 78766 3108 78818
rect 3052 78596 3108 78766
rect 3052 78530 3108 78540
rect 3276 75124 3332 79326
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 3500 78596 3556 78606
rect 3500 78502 3556 78540
rect 5852 78596 5908 78606
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 4396 76244 4452 76282
rect 4396 76178 4452 76188
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 3276 75058 3332 75068
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 3276 71652 3332 71662
rect 3276 71650 3444 71652
rect 3276 71598 3278 71650
rect 3330 71598 3444 71650
rect 3276 71596 3444 71598
rect 3276 71586 3332 71596
rect 3388 70980 3444 71596
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 3388 70914 3444 70924
rect 3388 70420 3444 70430
rect 3388 70326 3444 70364
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 3052 68626 3108 68638
rect 3052 68574 3054 68626
rect 3106 68574 3108 68626
rect 3052 68404 3108 68574
rect 3052 68338 3108 68348
rect 3612 68514 3668 68526
rect 3612 68462 3614 68514
rect 3666 68462 3668 68514
rect 3612 68404 3668 68462
rect 3612 68338 3668 68348
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 2940 67172 3220 67228
rect 1932 66164 1988 66174
rect 1820 66162 1988 66164
rect 1820 66110 1934 66162
rect 1986 66110 1988 66162
rect 1820 66108 1988 66110
rect 1820 65828 1876 66108
rect 1932 66098 1988 66108
rect 1820 65714 1876 65772
rect 1820 65662 1822 65714
rect 1874 65662 1876 65714
rect 1820 65650 1876 65662
rect 1820 64484 1876 64494
rect 1820 64482 1988 64484
rect 1820 64430 1822 64482
rect 1874 64430 1988 64482
rect 1820 64428 1988 64430
rect 1820 64418 1876 64428
rect 1932 64034 1988 64428
rect 1932 63982 1934 64034
rect 1986 63982 1988 64034
rect 1932 63364 1988 63982
rect 1932 63298 1988 63308
rect 1932 63028 1988 63038
rect 1820 63026 1988 63028
rect 1820 62974 1934 63026
rect 1986 62974 1988 63026
rect 1820 62972 1988 62974
rect 1820 62580 1876 62972
rect 1932 62962 1988 62972
rect 1820 62486 1876 62524
rect 3052 61684 3108 61694
rect 3052 61570 3108 61628
rect 3052 61518 3054 61570
rect 3106 61518 3108 61570
rect 3052 61506 3108 61518
rect 1932 61458 1988 61470
rect 1932 61406 1934 61458
rect 1986 61406 1988 61458
rect 1932 61348 1988 61406
rect 1932 61282 1988 61292
rect 1820 60676 1876 60686
rect 1820 60674 1988 60676
rect 1820 60622 1822 60674
rect 1874 60622 1988 60674
rect 1820 60620 1988 60622
rect 1820 60610 1876 60620
rect 1932 59892 1988 60620
rect 1932 59798 1988 59836
rect 1932 59332 1988 59342
rect 1820 59330 1988 59332
rect 1820 59278 1934 59330
rect 1986 59278 1988 59330
rect 1820 59276 1988 59278
rect 1820 58548 1876 59276
rect 1932 59266 1988 59276
rect 1820 58454 1876 58492
rect 3052 56866 3108 56878
rect 3052 56814 3054 56866
rect 3106 56814 3108 56866
rect 1932 56754 1988 56766
rect 1932 56702 1934 56754
rect 1986 56702 1988 56754
rect 1932 56644 1988 56702
rect 1932 56578 1988 56588
rect 3052 56644 3108 56814
rect 3052 56578 3108 56588
rect 1820 55074 1876 55086
rect 1820 55022 1822 55074
rect 1874 55022 1876 55074
rect 1820 54628 1876 55022
rect 1820 54562 1876 54572
rect 1932 52052 1988 52062
rect 1820 52050 1988 52052
rect 1820 51998 1934 52050
rect 1986 51998 1988 52050
rect 1820 51996 1988 51998
rect 1820 51716 1876 51996
rect 1932 51986 1988 51996
rect 1820 51602 1876 51660
rect 1820 51550 1822 51602
rect 1874 51550 1876 51602
rect 1820 51538 1876 51550
rect 1820 48802 1876 48814
rect 1820 48750 1822 48802
rect 1874 48750 1876 48802
rect 1820 48580 1876 48750
rect 1820 48514 1876 48524
rect 3164 47572 3220 67172
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 3276 66388 3332 66398
rect 3276 66294 3332 66332
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 3388 64148 3444 64158
rect 3276 63812 3332 63822
rect 3388 63812 3444 64092
rect 3276 63810 3444 63812
rect 3276 63758 3278 63810
rect 3330 63758 3444 63810
rect 3276 63756 3444 63758
rect 3276 63746 3332 63756
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 3276 63252 3332 63262
rect 5852 63252 5908 78540
rect 7532 69748 7588 116510
rect 9884 116564 9940 116574
rect 10108 116564 10164 119200
rect 9884 116562 10500 116564
rect 9884 116510 9886 116562
rect 9938 116510 10500 116562
rect 9884 116508 10500 116510
rect 9884 116498 9940 116508
rect 10444 116338 10500 116508
rect 10444 116286 10446 116338
rect 10498 116286 10500 116338
rect 10444 116274 10500 116286
rect 10668 115778 10724 115790
rect 10668 115726 10670 115778
rect 10722 115726 10724 115778
rect 10332 115666 10388 115678
rect 10332 115614 10334 115666
rect 10386 115614 10388 115666
rect 9772 115556 9828 115566
rect 9772 115462 9828 115500
rect 10332 115556 10388 115614
rect 10668 115668 10724 115726
rect 11228 115668 11284 115678
rect 10668 115666 11284 115668
rect 10668 115614 11230 115666
rect 11282 115614 11284 115666
rect 10668 115612 11284 115614
rect 11228 115602 11284 115612
rect 10332 115490 10388 115500
rect 11340 115556 11396 115566
rect 11564 115556 11620 119200
rect 11788 116564 11844 116574
rect 11788 116470 11844 116508
rect 12796 116562 12852 119200
rect 16044 117460 16100 119200
rect 12796 116510 12798 116562
rect 12850 116510 12852 116562
rect 12796 115780 12852 116510
rect 15708 117404 16100 117460
rect 15708 116452 15764 117404
rect 16716 116564 16772 116574
rect 16716 116562 16884 116564
rect 16716 116510 16718 116562
rect 16770 116510 16884 116562
rect 16716 116508 16884 116510
rect 16716 116498 16772 116508
rect 15708 116338 15764 116396
rect 15708 116286 15710 116338
rect 15762 116286 15764 116338
rect 15708 116274 15764 116286
rect 13132 115780 13188 115790
rect 12796 115778 13188 115780
rect 12796 115726 13134 115778
rect 13186 115726 13188 115778
rect 12796 115724 13188 115726
rect 13132 115714 13188 115724
rect 12348 115668 12404 115678
rect 11900 115556 11956 115566
rect 11564 115554 11956 115556
rect 11564 115502 11902 115554
rect 11954 115502 11956 115554
rect 11564 115500 11956 115502
rect 11340 114994 11396 115500
rect 11900 115490 11956 115500
rect 12348 114996 12404 115612
rect 11340 114942 11342 114994
rect 11394 114942 11396 114994
rect 11340 114930 11396 114942
rect 11900 114994 12404 114996
rect 11900 114942 12350 114994
rect 12402 114942 12404 114994
rect 11900 114940 12404 114942
rect 11900 114882 11956 114940
rect 12348 114930 12404 114940
rect 14252 115554 14308 115566
rect 14252 115502 14254 115554
rect 14306 115502 14308 115554
rect 11900 114830 11902 114882
rect 11954 114830 11956 114882
rect 11900 114660 11956 114830
rect 11900 114594 11956 114604
rect 7532 69682 7588 69692
rect 9212 113988 9268 113998
rect 3276 63250 3556 63252
rect 3276 63198 3278 63250
rect 3330 63198 3556 63250
rect 3276 63196 3556 63198
rect 3276 63186 3332 63196
rect 3388 60228 3444 60238
rect 3276 60172 3388 60228
rect 3276 60114 3332 60172
rect 3388 60162 3444 60172
rect 3276 60062 3278 60114
rect 3330 60062 3332 60114
rect 3276 60050 3332 60062
rect 3276 59108 3332 59118
rect 3276 59014 3332 59052
rect 3500 58212 3556 63196
rect 5852 63186 5908 63196
rect 6748 68516 6804 68526
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 3612 61684 3668 61694
rect 3612 61590 3668 61628
rect 6748 61684 6804 68460
rect 6748 61618 6804 61628
rect 5852 60900 5908 60910
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 5852 60228 5908 60844
rect 5852 60162 5908 60172
rect 5852 59444 5908 59454
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 3500 58146 3556 58156
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 3500 56644 3556 56654
rect 3500 56550 3556 56588
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3276 52274 3332 52286
rect 3276 52222 3278 52274
rect 3330 52222 3332 52274
rect 3276 52052 3332 52222
rect 3388 52052 3444 52062
rect 3276 51996 3388 52052
rect 3388 51986 3444 51996
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 3276 47572 3332 47582
rect 2604 47570 3332 47572
rect 2604 47518 3278 47570
rect 3330 47518 3332 47570
rect 2604 47516 3332 47518
rect 2604 47458 2660 47516
rect 2604 47406 2606 47458
rect 2658 47406 2660 47458
rect 2604 47394 2660 47406
rect 2828 47234 2884 47246
rect 2828 47182 2830 47234
rect 2882 47182 2884 47234
rect 2828 46674 2884 47182
rect 2828 46622 2830 46674
rect 2882 46622 2884 46674
rect 2828 46610 2884 46622
rect 1932 46564 1988 46574
rect 1932 46470 1988 46508
rect 3052 45890 3108 45902
rect 3052 45838 3054 45890
rect 3106 45838 3108 45890
rect 1932 45778 1988 45790
rect 1932 45726 1934 45778
rect 1986 45726 1988 45778
rect 1932 45220 1988 45726
rect 3052 45668 3108 45838
rect 3052 45602 3108 45612
rect 1932 45154 1988 45164
rect 1932 41076 1988 41086
rect 1708 41074 1988 41076
rect 1708 41022 1934 41074
rect 1986 41022 1988 41074
rect 1708 41020 1988 41022
rect 1708 40516 1764 41020
rect 1932 41010 1988 41020
rect 1708 40422 1764 40460
rect 3052 39620 3108 39630
rect 3052 39526 3108 39564
rect 1932 39506 1988 39518
rect 1932 39454 1934 39506
rect 1986 39454 1988 39506
rect 1932 39172 1988 39454
rect 1932 39106 1988 39116
rect 3052 38050 3108 38062
rect 3052 37998 3054 38050
rect 3106 37998 3108 38050
rect 1932 37938 1988 37950
rect 1932 37886 1934 37938
rect 1986 37886 1988 37938
rect 1932 37828 1988 37886
rect 1932 37762 1988 37772
rect 3052 37828 3108 37998
rect 3052 37762 3108 37772
rect 1932 37378 1988 37390
rect 1932 37326 1934 37378
rect 1986 37326 1988 37378
rect 1932 37156 1988 37326
rect 1820 35924 1876 35934
rect 1932 35924 1988 37100
rect 1820 35922 1988 35924
rect 1820 35870 1822 35922
rect 1874 35870 1988 35922
rect 1820 35868 1988 35870
rect 2156 36370 2212 36382
rect 2156 36318 2158 36370
rect 2210 36318 2212 36370
rect 1820 35858 1876 35868
rect 2156 35812 2212 36318
rect 2156 35718 2212 35756
rect 1932 34802 1988 34814
rect 1932 34750 1934 34802
rect 1986 34750 1988 34802
rect 1932 34468 1988 34750
rect 1820 34412 1932 34468
rect 1820 33458 1876 34412
rect 1932 34402 1988 34412
rect 3052 34130 3108 34142
rect 3052 34078 3054 34130
rect 3106 34078 3108 34130
rect 1932 34018 1988 34030
rect 1932 33966 1934 34018
rect 1986 33966 1988 34018
rect 1932 33796 1988 33966
rect 3052 34020 3108 34078
rect 3052 33954 3108 33964
rect 1932 33730 1988 33740
rect 1820 33406 1822 33458
rect 1874 33406 1876 33458
rect 1820 33394 1876 33406
rect 1932 32674 1988 32686
rect 1932 32622 1934 32674
rect 1986 32622 1988 32674
rect 1932 32228 1988 32622
rect 1932 31948 1988 32172
rect 1820 31892 1988 31948
rect 1820 31890 1876 31892
rect 1820 31838 1822 31890
rect 1874 31838 1876 31890
rect 1820 31826 1876 31838
rect 1932 30100 1988 30110
rect 1820 30098 1988 30100
rect 1820 30046 1934 30098
rect 1986 30046 1988 30098
rect 1820 30044 1988 30046
rect 1820 29652 1876 30044
rect 1932 30034 1988 30044
rect 1820 29558 1876 29596
rect 1932 26964 1988 26974
rect 1708 26962 1988 26964
rect 1708 26910 1934 26962
rect 1986 26910 1988 26962
rect 1708 26908 1988 26910
rect 1708 26404 1764 26908
rect 1932 26898 1988 26908
rect 1708 26310 1764 26348
rect 2156 26178 2212 26190
rect 2156 26126 2158 26178
rect 2210 26126 2212 26178
rect 1932 25396 1988 25406
rect 2156 25396 2212 26126
rect 1932 25394 2212 25396
rect 1932 25342 1934 25394
rect 1986 25342 2212 25394
rect 1932 25340 2212 25342
rect 1932 25060 1988 25340
rect 1932 24994 1988 25004
rect 3052 24722 3108 24734
rect 3052 24670 3054 24722
rect 3106 24670 3108 24722
rect 1932 24610 1988 24622
rect 1932 24558 1934 24610
rect 1986 24558 1988 24610
rect 1932 24388 1988 24558
rect 3052 24612 3108 24670
rect 3052 24546 3108 24556
rect 1932 24322 1988 24332
rect 3052 23154 3108 23166
rect 3052 23102 3054 23154
rect 3106 23102 3108 23154
rect 1932 23044 1988 23054
rect 1932 22950 1988 22988
rect 3052 23044 3108 23102
rect 3052 22978 3108 22988
rect 1932 22260 1988 22270
rect 1820 22258 1988 22260
rect 1820 22206 1934 22258
rect 1986 22206 1988 22258
rect 1820 22204 1988 22206
rect 1820 21476 1876 22204
rect 1932 22194 1988 22204
rect 3052 21586 3108 21598
rect 3052 21534 3054 21586
rect 3106 21534 3108 21586
rect 1820 20914 1876 21420
rect 1932 21474 1988 21486
rect 1932 21422 1934 21474
rect 1986 21422 1988 21474
rect 1932 21028 1988 21422
rect 3052 21364 3108 21534
rect 3052 21298 3108 21308
rect 1932 20962 1988 20972
rect 1820 20862 1822 20914
rect 1874 20862 1876 20914
rect 1820 20850 1876 20862
rect 1820 18562 1876 18574
rect 1820 18510 1822 18562
rect 1874 18510 1876 18562
rect 1820 18340 1876 18510
rect 1820 18274 1876 18284
rect 1820 17442 1876 17454
rect 1820 17390 1822 17442
rect 1874 17390 1876 17442
rect 1820 16996 1876 17390
rect 1820 16930 1876 16940
rect 3052 16884 3108 16894
rect 3052 16790 3108 16828
rect 1932 16770 1988 16782
rect 1932 16718 1934 16770
rect 1986 16718 1988 16770
rect 1932 16324 1988 16718
rect 1932 16258 1988 16268
rect 2828 12178 2884 12190
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 1932 12066 1988 12078
rect 1932 12014 1934 12066
rect 1986 12014 1988 12066
rect 1932 11620 1988 12014
rect 1932 11554 1988 11564
rect 2604 11394 2660 11406
rect 2604 11342 2606 11394
rect 2658 11342 2660 11394
rect 2604 11060 2660 11342
rect 2828 11282 2884 12126
rect 2828 11230 2830 11282
rect 2882 11230 2884 11282
rect 2828 11218 2884 11230
rect 3164 11508 3220 47516
rect 3276 47506 3332 47516
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 3500 45668 3556 45678
rect 3500 45574 3556 45612
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 3276 41300 3332 41310
rect 3276 41206 3332 41244
rect 3612 41188 3668 41198
rect 3612 39730 3668 41132
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 3612 39678 3614 39730
rect 3666 39678 3668 39730
rect 3612 39620 3668 39678
rect 3612 39554 3668 39564
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 3388 37940 3444 37950
rect 3276 37156 3332 37166
rect 3388 37156 3444 37884
rect 3500 37828 3556 37838
rect 3500 37734 3556 37772
rect 3276 37154 3444 37156
rect 3276 37102 3278 37154
rect 3330 37102 3444 37154
rect 3276 37100 3444 37102
rect 3276 37090 3332 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 3276 36596 3332 36606
rect 3276 36502 3332 36540
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3388 35140 3444 35150
rect 3276 35028 3332 35038
rect 3388 35028 3444 35084
rect 3276 35026 3444 35028
rect 3276 34974 3278 35026
rect 3330 34974 3444 35026
rect 3276 34972 3444 34974
rect 3276 34962 3332 34972
rect 3612 34020 3668 34030
rect 3612 33926 3668 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 3276 32452 3332 32462
rect 3276 32358 3332 32396
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 3276 30322 3332 30334
rect 3276 30270 3278 30322
rect 3330 30270 3332 30322
rect 3276 30212 3332 30270
rect 3388 30212 3444 30222
rect 3276 30156 3388 30212
rect 3388 30146 3444 30156
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3388 27300 3444 27310
rect 3276 27244 3388 27300
rect 3276 27186 3332 27244
rect 3388 27234 3444 27244
rect 3276 27134 3278 27186
rect 3330 27134 3332 27186
rect 3276 27122 3332 27134
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3388 25732 3444 25742
rect 3276 25676 3388 25732
rect 3276 25618 3332 25676
rect 3388 25666 3444 25676
rect 5852 25732 5908 59388
rect 9212 57764 9268 113932
rect 9212 57698 9268 57708
rect 10892 70980 10948 70990
rect 7532 49588 7588 49598
rect 7532 27300 7588 49532
rect 8428 46788 8484 46798
rect 8428 37940 8484 46732
rect 10892 43428 10948 70924
rect 10892 43362 10948 43372
rect 12908 66164 12964 66174
rect 10556 42868 10612 42878
rect 8428 37874 8484 37884
rect 8764 39732 8820 39742
rect 8764 35140 8820 39676
rect 8764 35074 8820 35084
rect 7532 27234 7588 27244
rect 5852 25666 5908 25676
rect 9660 27076 9716 27086
rect 3276 25566 3278 25618
rect 3330 25566 3332 25618
rect 3276 25554 3332 25566
rect 3500 24612 3556 24622
rect 3500 24518 3556 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 3500 23044 3556 23054
rect 3500 22950 3556 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4396 22148 4452 22158
rect 4396 22054 4452 22092
rect 3612 21474 3668 21486
rect 3612 21422 3614 21474
rect 3666 21422 3668 21474
rect 3612 21364 3668 21422
rect 3612 21298 3668 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5628 19796 5684 19806
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3500 16884 3556 16894
rect 3500 16790 3556 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 3276 11508 3332 11518
rect 3164 11506 3332 11508
rect 3164 11454 3278 11506
rect 3330 11454 3332 11506
rect 3164 11452 3332 11454
rect 3164 11060 3220 11452
rect 3276 11442 3332 11452
rect 2604 11004 3220 11060
rect 3052 10610 3108 10622
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 1932 10498 1988 10510
rect 1932 10446 1934 10498
rect 1986 10446 1988 10498
rect 1932 10276 1988 10446
rect 3052 10500 3108 10558
rect 3052 10434 3108 10444
rect 1932 10210 1988 10220
rect 1820 7586 1876 7598
rect 1820 7534 1822 7586
rect 1874 7534 1876 7586
rect 1820 6916 1876 7534
rect 1820 6850 1876 6860
rect 2380 7362 2436 7374
rect 2380 7310 2382 7362
rect 2434 7310 2436 7362
rect 1932 6580 1988 6590
rect 1932 6578 2100 6580
rect 1932 6526 1934 6578
rect 1986 6526 2100 6578
rect 1932 6524 2100 6526
rect 1932 6514 1988 6524
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5572 1988 5742
rect 1932 5506 1988 5516
rect 1932 5012 1988 5022
rect 1820 5010 1988 5012
rect 1820 4958 1934 5010
rect 1986 4958 1988 5010
rect 1820 4956 1988 4958
rect 812 4452 868 4462
rect 140 3668 196 3678
rect 140 800 196 3612
rect 812 800 868 4396
rect 1820 4228 1876 4956
rect 1932 4946 1988 4956
rect 1932 4452 1988 4462
rect 1932 4358 1988 4396
rect 1820 4162 1876 4172
rect 2044 3668 2100 6524
rect 2380 4452 2436 7310
rect 3052 6690 3108 6702
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6468 3108 6638
rect 3052 6402 3108 6412
rect 3052 5908 3108 5918
rect 3052 5814 3108 5852
rect 2828 5124 2884 5134
rect 2380 4386 2436 4396
rect 2492 5122 2884 5124
rect 2492 5070 2830 5122
rect 2882 5070 2884 5122
rect 2492 5068 2884 5070
rect 2044 3602 2100 3612
rect 2156 4228 2212 4238
rect 2044 3444 2100 3454
rect 2044 3350 2100 3388
rect 2156 800 2212 4172
rect 2492 3330 2548 5068
rect 2828 5058 2884 5068
rect 2828 4340 2884 4350
rect 2828 3554 2884 4284
rect 3164 4340 3220 11004
rect 3500 10500 3556 10510
rect 3500 10406 3556 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 3612 6468 3668 6478
rect 3612 6374 3668 6412
rect 3500 5908 3556 5918
rect 3500 5814 3556 5852
rect 3836 5796 3892 5806
rect 3724 5010 3780 5022
rect 3724 4958 3726 5010
rect 3778 4958 3780 5010
rect 3164 4274 3220 4284
rect 3388 4452 3444 4462
rect 3276 4228 3332 4238
rect 3388 4228 3444 4396
rect 3276 4226 3444 4228
rect 3276 4174 3278 4226
rect 3330 4174 3444 4226
rect 3276 4172 3444 4174
rect 3276 4162 3332 4172
rect 2828 3502 2830 3554
rect 2882 3502 2884 3554
rect 2828 3444 2884 3502
rect 3724 3556 3780 4958
rect 3724 3490 3780 3500
rect 2828 3378 2884 3388
rect 3500 3444 3556 3454
rect 2492 3278 2494 3330
rect 2546 3278 2548 3330
rect 2492 3266 2548 3278
rect 3500 2212 3556 3388
rect 3836 3444 3892 5740
rect 5180 5796 5236 5806
rect 5180 5702 5236 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4956 5236 5012 5246
rect 4844 5124 4900 5134
rect 4844 5030 4900 5068
rect 4956 4338 5012 5180
rect 5628 5234 5684 19740
rect 5628 5182 5630 5234
rect 5682 5182 5684 5234
rect 5628 5124 5684 5182
rect 6076 5236 6132 5246
rect 6076 5142 6132 5180
rect 5628 4450 5684 5068
rect 6524 5124 6580 5134
rect 6524 4562 6580 5068
rect 9660 4564 9716 27020
rect 6524 4510 6526 4562
rect 6578 4510 6580 4562
rect 6524 4498 6580 4510
rect 8876 4562 9716 4564
rect 8876 4510 9662 4562
rect 9714 4510 9716 4562
rect 8876 4508 9716 4510
rect 5628 4398 5630 4450
rect 5682 4398 5684 4450
rect 5628 4386 5684 4398
rect 5964 4450 6020 4462
rect 5964 4398 5966 4450
rect 6018 4398 6020 4450
rect 4956 4286 4958 4338
rect 5010 4286 5012 4338
rect 4956 4274 5012 4286
rect 3948 4228 4004 4238
rect 3948 4134 4004 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4956 3668 5012 3678
rect 4956 3574 5012 3612
rect 5964 3554 6020 4398
rect 8204 4338 8260 4350
rect 8204 4286 8206 4338
rect 8258 4286 8260 4338
rect 7084 4226 7140 4238
rect 7084 4174 7086 4226
rect 7138 4174 7140 4226
rect 5964 3502 5966 3554
rect 6018 3502 6020 3554
rect 5964 3490 6020 3502
rect 6412 3666 6468 3678
rect 6412 3614 6414 3666
rect 6466 3614 6468 3666
rect 6412 3444 6468 3614
rect 3836 3442 4004 3444
rect 3836 3390 3838 3442
rect 3890 3390 4004 3442
rect 3836 3388 4004 3390
rect 3836 3378 3892 3388
rect 3500 2146 3556 2156
rect 3948 800 4004 3388
rect 6412 3378 6468 3388
rect 7084 868 7140 4174
rect 8204 4228 8260 4286
rect 8204 4162 8260 4172
rect 8764 4228 8820 4238
rect 8764 4134 8820 4172
rect 8876 4004 8932 4508
rect 9660 4498 9716 4508
rect 10556 4562 10612 42812
rect 12348 31220 12404 31230
rect 12348 23044 12404 31164
rect 12348 22978 12404 22988
rect 10556 4510 10558 4562
rect 10610 4510 10612 4562
rect 8764 3948 8932 4004
rect 6860 812 7140 868
rect 7980 3666 8036 3678
rect 7980 3614 7982 3666
rect 8034 3614 8036 3666
rect 6860 800 6916 812
rect -56 728 196 800
rect 616 728 868 800
rect 1960 728 2212 800
rect -56 200 168 728
rect 616 200 840 728
rect 1960 200 2184 728
rect 3304 200 3528 800
rect 3948 728 4200 800
rect 3976 200 4200 728
rect 5320 200 5544 800
rect 6664 728 6916 800
rect 7980 800 8036 3614
rect 8764 3554 8820 3948
rect 8764 3502 8766 3554
rect 8818 3502 8820 3554
rect 8764 3490 8820 3502
rect 10556 3556 10612 4510
rect 11228 4564 11284 4574
rect 11228 4340 11284 4508
rect 11900 4564 11956 4574
rect 11900 4470 11956 4508
rect 11452 4452 11508 4462
rect 11452 4450 11620 4452
rect 11452 4398 11454 4450
rect 11506 4398 11620 4450
rect 11452 4396 11620 4398
rect 11452 4386 11508 4396
rect 11228 4208 11284 4284
rect 11452 3668 11508 3678
rect 10668 3556 10724 3566
rect 10556 3554 10724 3556
rect 10556 3502 10670 3554
rect 10722 3502 10724 3554
rect 10556 3500 10724 3502
rect 10668 3490 10724 3500
rect 8876 3444 8932 3454
rect 8876 800 8932 3388
rect 9772 3444 9828 3454
rect 9772 3350 9828 3388
rect 11452 800 11508 3612
rect 11564 3554 11620 4396
rect 12908 3780 12964 66108
rect 14252 64708 14308 115502
rect 15932 97748 15988 97758
rect 15932 68068 15988 97692
rect 16828 69972 16884 116508
rect 17388 116452 17444 116462
rect 17388 116358 17444 116396
rect 18956 116340 19012 119200
rect 20972 116564 21028 116574
rect 19068 116340 19124 116350
rect 18956 116338 19124 116340
rect 18956 116286 19070 116338
rect 19122 116286 19124 116338
rect 18956 116284 19124 116286
rect 19068 116274 19124 116284
rect 19836 116060 20100 116070
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 19836 115994 20100 116004
rect 19836 114492 20100 114502
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 19836 114426 20100 114436
rect 19836 112924 20100 112934
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 19836 112858 20100 112868
rect 19836 111356 20100 111366
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 19836 111290 20100 111300
rect 19836 109788 20100 109798
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 19836 109722 20100 109732
rect 19836 108220 20100 108230
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 19836 108154 20100 108164
rect 19836 106652 20100 106662
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 19836 106586 20100 106596
rect 19836 105084 20100 105094
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 19836 105018 20100 105028
rect 19836 103516 20100 103526
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 19836 103450 20100 103460
rect 19836 101948 20100 101958
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 19836 101882 20100 101892
rect 19836 100380 20100 100390
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 19836 100314 20100 100324
rect 19836 98812 20100 98822
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 19836 98746 20100 98756
rect 19836 97244 20100 97254
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 19836 97178 20100 97188
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 16828 69906 16884 69916
rect 17612 69748 17668 69758
rect 15932 68002 15988 68012
rect 16156 68404 16212 68414
rect 14252 64642 14308 64652
rect 14252 48356 14308 48366
rect 13580 16884 13636 16894
rect 13580 15204 13636 16828
rect 13580 15138 13636 15148
rect 14252 4452 14308 48300
rect 16156 47684 16212 68348
rect 17612 56868 17668 69692
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 20972 63364 21028 116508
rect 21980 116564 22036 116574
rect 22092 116564 22148 119200
rect 21980 116562 22148 116564
rect 21980 116510 21982 116562
rect 22034 116510 22148 116562
rect 21980 116508 22148 116510
rect 21980 116498 22036 116508
rect 22092 116340 22148 116508
rect 23884 116564 23940 116574
rect 24332 116564 24388 119200
rect 23884 116562 24164 116564
rect 23884 116510 23886 116562
rect 23938 116510 24164 116562
rect 23884 116508 24164 116510
rect 23884 116498 23940 116508
rect 23548 116452 23604 116462
rect 22540 116340 22596 116350
rect 22092 116338 22596 116340
rect 22092 116286 22542 116338
rect 22594 116286 22596 116338
rect 22092 116284 22596 116286
rect 22540 116274 22596 116284
rect 22764 115892 22820 115902
rect 22764 115798 22820 115836
rect 23548 115890 23604 116396
rect 23548 115838 23550 115890
rect 23602 115838 23604 115890
rect 23548 115826 23604 115838
rect 24108 115892 24164 116508
rect 24332 116498 24388 116508
rect 26012 116564 26068 116574
rect 26012 116470 26068 116508
rect 25340 116452 25396 116462
rect 25340 116358 25396 116396
rect 24108 115798 24164 115836
rect 28700 115892 28756 115902
rect 28812 115892 28868 119200
rect 31388 116340 31444 116350
rect 31500 116340 31556 119200
rect 32172 117460 32228 119200
rect 31388 116338 31500 116340
rect 31388 116286 31390 116338
rect 31442 116286 31500 116338
rect 31388 116284 31500 116286
rect 31388 116274 31444 116284
rect 31500 116208 31556 116284
rect 32060 117404 32228 117460
rect 28700 115890 28868 115892
rect 28700 115838 28702 115890
rect 28754 115838 28868 115890
rect 28700 115836 28868 115838
rect 28700 115826 28756 115836
rect 28812 115780 28868 115836
rect 29260 115780 29316 115790
rect 28812 115778 29316 115780
rect 28812 115726 29262 115778
rect 29314 115726 29316 115778
rect 28812 115724 29316 115726
rect 29260 115714 29316 115724
rect 23324 115668 23380 115678
rect 23324 114660 23380 115612
rect 24668 115554 24724 115566
rect 24668 115502 24670 115554
rect 24722 115502 24724 115554
rect 23324 114594 23380 114604
rect 23772 114660 23828 114670
rect 23772 114566 23828 114604
rect 24668 114660 24724 115502
rect 24668 114594 24724 114604
rect 30380 115554 30436 115566
rect 30380 115502 30382 115554
rect 30434 115502 30436 115554
rect 29372 111860 29428 111870
rect 20972 63298 21028 63308
rect 22652 102452 22708 102462
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 22652 62356 22708 102396
rect 22652 62290 22708 62300
rect 24332 88340 24388 88350
rect 24332 61348 24388 88284
rect 24332 61282 24388 61292
rect 26012 76244 26068 76254
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 20972 60004 21028 60014
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 17612 56802 17668 56812
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 16156 47618 16212 47628
rect 17612 51268 17668 51278
rect 15932 42532 15988 42542
rect 15932 30212 15988 42476
rect 15932 30146 15988 30156
rect 17612 24612 17668 51212
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 17612 24546 17668 24556
rect 17836 23940 17892 23950
rect 14252 4386 14308 4396
rect 15372 9268 15428 9278
rect 15372 4562 15428 9212
rect 17836 5908 17892 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 17836 5842 17892 5852
rect 19628 12740 19684 12750
rect 15372 4510 15374 4562
rect 15426 4510 15428 4562
rect 14924 4340 14980 4350
rect 15372 4340 15428 4510
rect 14924 4338 15428 4340
rect 14924 4286 14926 4338
rect 14978 4286 15428 4338
rect 14924 4284 15428 4286
rect 18508 4450 18564 4462
rect 18508 4398 18510 4450
rect 18562 4398 18564 4450
rect 14924 4274 14980 4284
rect 13804 4228 13860 4238
rect 12908 3714 12964 3724
rect 13580 4226 13860 4228
rect 13580 4174 13806 4226
rect 13858 4174 13860 4226
rect 13580 4172 13860 4174
rect 12236 3668 12292 3678
rect 12236 3574 12292 3612
rect 11564 3502 11566 3554
rect 11618 3502 11620 3554
rect 11564 3490 11620 3502
rect 13580 800 13636 4172
rect 13804 4162 13860 4172
rect 17948 4228 18004 4238
rect 18508 4228 18564 4398
rect 17948 4226 18564 4228
rect 17948 4174 17950 4226
rect 18002 4174 18564 4226
rect 17948 4172 18564 4174
rect 19628 4226 19684 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20972 5124 21028 59948
rect 26012 59332 26068 76188
rect 26012 59266 26068 59276
rect 26012 57428 26068 57438
rect 22652 56756 22708 56766
rect 22652 41300 22708 56700
rect 22652 41234 22708 41244
rect 24332 55076 24388 55086
rect 20972 5058 21028 5068
rect 22652 39844 22708 39854
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4174 19630 4226
rect 19682 4174 19684 4226
rect 17948 4162 18004 4172
rect 16492 3668 16548 3678
rect 16492 3574 16548 3612
rect 14588 3444 14644 3454
rect 15148 3444 15204 3454
rect 14588 3442 15204 3444
rect 14588 3390 14590 3442
rect 14642 3390 15150 3442
rect 15202 3390 15204 3442
rect 14588 3388 15204 3390
rect 14588 3378 14644 3388
rect 7980 728 8232 800
rect 6664 200 6888 728
rect 8008 200 8232 728
rect 8680 728 8932 800
rect 8680 200 8904 728
rect 10024 200 10248 800
rect 11368 200 11592 800
rect 12040 200 12264 800
rect 13384 728 13636 800
rect 14700 800 14756 3388
rect 15148 3378 15204 3388
rect 18060 800 18116 4172
rect 19628 4162 19684 4174
rect 21196 4226 21252 4238
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 19628 3892 19684 3902
rect 19628 3442 19684 3836
rect 20636 3780 20692 3790
rect 20636 3666 20692 3724
rect 20636 3614 20638 3666
rect 20690 3614 20692 3666
rect 20636 3602 20692 3614
rect 19628 3390 19630 3442
rect 19682 3390 19684 3442
rect 19628 800 19684 3390
rect 20972 3444 21028 3454
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20972 800 21028 3388
rect 21196 3444 21252 4174
rect 21532 4226 21588 4238
rect 21532 4174 21534 4226
rect 21586 4174 21588 4226
rect 21532 3892 21588 4174
rect 21532 3826 21588 3836
rect 22652 3666 22708 39788
rect 22652 3614 22654 3666
rect 22706 3614 22708 3666
rect 22652 3602 22708 3614
rect 24332 3668 24388 55020
rect 26012 22148 26068 57372
rect 29372 51604 29428 111804
rect 30380 53508 30436 115502
rect 32060 115554 32116 117404
rect 33740 117124 33796 119200
rect 33740 117068 34020 117124
rect 32060 115502 32062 115554
rect 32114 115502 32116 115554
rect 32060 115490 32116 115502
rect 32172 116562 32228 116574
rect 32172 116510 32174 116562
rect 32226 116510 32228 116562
rect 32172 101780 32228 116510
rect 33068 116340 33124 116350
rect 33068 116246 33124 116284
rect 32844 115666 32900 115678
rect 32844 115614 32846 115666
rect 32898 115614 32900 115666
rect 32844 115556 32900 115614
rect 32844 115490 32900 115500
rect 33628 115556 33684 115566
rect 33628 115462 33684 115500
rect 33964 114994 34020 117068
rect 35084 115780 35140 119200
rect 35532 119200 35784 119336
rect 36904 119200 37128 119800
rect 38248 119336 38472 119800
rect 38220 119200 38472 119336
rect 39592 119336 39816 119800
rect 39592 119200 39844 119336
rect 40264 119200 40488 119800
rect 41608 119336 41832 119800
rect 42952 119336 43176 119800
rect 41608 119200 41860 119336
rect 42952 119200 43204 119336
rect 43624 119200 43848 119800
rect 44968 119200 45192 119800
rect 46312 119336 46536 119800
rect 47656 119336 47880 119800
rect 46312 119200 46564 119336
rect 35196 116844 35460 116854
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35196 116778 35460 116788
rect 35532 116564 35588 119200
rect 35196 116340 35252 116350
rect 35532 116340 35588 116508
rect 35196 116338 35588 116340
rect 35196 116286 35198 116338
rect 35250 116286 35588 116338
rect 35196 116284 35588 116286
rect 36316 116562 36372 116574
rect 36316 116510 36318 116562
rect 36370 116510 36372 116562
rect 35196 116274 35252 116284
rect 36316 116004 36372 116510
rect 36316 115938 36372 115948
rect 36988 116562 37044 119200
rect 36988 116510 36990 116562
rect 37042 116510 37044 116562
rect 35308 115780 35364 115790
rect 35084 115778 35364 115780
rect 35084 115726 35310 115778
rect 35362 115726 35364 115778
rect 35084 115724 35364 115726
rect 36988 115780 37044 116510
rect 37436 116564 37492 116574
rect 37436 116470 37492 116508
rect 38108 116564 38164 116574
rect 38220 116564 38276 119200
rect 39788 117122 39844 119200
rect 39788 117070 39790 117122
rect 39842 117070 39844 117122
rect 39788 117058 39844 117070
rect 41132 117122 41188 117134
rect 41132 117070 41134 117122
rect 41186 117070 41188 117122
rect 38108 116562 38276 116564
rect 38108 116510 38110 116562
rect 38162 116510 38276 116562
rect 38108 116508 38276 116510
rect 38108 116498 38164 116508
rect 38220 116340 38276 116508
rect 39788 116562 39844 116574
rect 39788 116510 39790 116562
rect 39842 116510 39844 116562
rect 38668 116340 38724 116350
rect 38220 116338 38724 116340
rect 38220 116286 38670 116338
rect 38722 116286 38724 116338
rect 38220 116284 38724 116286
rect 38668 116274 38724 116284
rect 37324 115780 37380 115790
rect 36988 115778 37380 115780
rect 36988 115726 37326 115778
rect 37378 115726 37380 115778
rect 36988 115724 37380 115726
rect 35308 115714 35364 115724
rect 37324 115714 37380 115724
rect 36428 115668 36484 115678
rect 36428 115666 36708 115668
rect 36428 115614 36430 115666
rect 36482 115614 36708 115666
rect 36428 115612 36708 115614
rect 36428 115602 36484 115612
rect 35196 115276 35460 115286
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35196 115210 35460 115220
rect 33964 114942 33966 114994
rect 34018 114942 34020 114994
rect 33964 114930 34020 114942
rect 36652 114994 36708 115612
rect 36652 114942 36654 114994
rect 36706 114942 36708 114994
rect 34860 114882 34916 114894
rect 34860 114830 34862 114882
rect 34914 114830 34916 114882
rect 33964 114660 34020 114670
rect 32172 101714 32228 101724
rect 32732 104580 32788 104590
rect 32732 66500 32788 104524
rect 32732 66434 32788 66444
rect 32172 66388 32228 66398
rect 32172 59668 32228 66332
rect 32172 59602 32228 59612
rect 33516 59108 33572 59118
rect 33516 55972 33572 59052
rect 33516 55906 33572 55916
rect 30380 53442 30436 53452
rect 33516 54404 33572 54414
rect 29372 51538 29428 51548
rect 31052 52164 31108 52174
rect 27020 48916 27076 48926
rect 26012 22082 26068 22092
rect 26124 23716 26180 23726
rect 26124 10500 26180 23660
rect 26124 10434 26180 10444
rect 25228 5124 25284 5134
rect 24332 3602 24388 3612
rect 25004 5122 25284 5124
rect 25004 5070 25230 5122
rect 25282 5070 25284 5122
rect 25004 5068 25284 5070
rect 21196 3378 21252 3388
rect 21532 3444 21588 3454
rect 21532 3350 21588 3388
rect 24668 3444 24724 3454
rect 24332 812 24500 868
rect 24332 800 24388 812
rect 14700 728 14952 800
rect 13384 200 13608 728
rect 14728 200 14952 728
rect 16072 200 16296 800
rect 16744 200 16968 800
rect 18060 728 18312 800
rect 18088 200 18312 728
rect 19432 728 19684 800
rect 20776 728 21028 800
rect 19432 200 19656 728
rect 20776 200 21000 728
rect 21448 200 21672 800
rect 22792 200 23016 800
rect 24136 728 24388 800
rect 24444 756 24500 812
rect 24668 756 24724 3388
rect 25004 800 25060 5068
rect 25228 5058 25284 5068
rect 26348 5124 26404 5134
rect 26348 5030 26404 5068
rect 26908 5124 26964 5134
rect 26908 5030 26964 5068
rect 26572 4228 26628 4238
rect 26348 4226 26628 4228
rect 26348 4174 26574 4226
rect 26626 4174 26628 4226
rect 26348 4172 26628 4174
rect 25452 3444 25508 3454
rect 25452 3350 25508 3388
rect 26348 800 26404 4172
rect 26572 4162 26628 4172
rect 26796 3668 26852 3678
rect 27020 3668 27076 48860
rect 29372 44884 29428 44894
rect 29372 12740 29428 44828
rect 29372 12674 29428 12684
rect 29484 26964 29540 26974
rect 29484 6468 29540 26908
rect 29484 6402 29540 6412
rect 28140 5236 28196 5246
rect 28140 4562 28196 5180
rect 28140 4510 28142 4562
rect 28194 4510 28196 4562
rect 27692 4340 27748 4350
rect 28140 4340 28196 4510
rect 27692 4338 28196 4340
rect 27692 4286 27694 4338
rect 27746 4286 28196 4338
rect 27692 4284 28196 4286
rect 27692 4274 27748 4284
rect 26796 3666 27076 3668
rect 26796 3614 26798 3666
rect 26850 3614 27076 3666
rect 26796 3612 27076 3614
rect 31052 3666 31108 52108
rect 33516 52164 33572 54348
rect 33964 53170 34020 114604
rect 34860 114660 34916 114830
rect 34860 114594 34916 114604
rect 35532 114660 35588 114670
rect 35532 114566 35588 114604
rect 35196 113708 35460 113718
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35196 113642 35460 113652
rect 35196 112140 35460 112150
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35196 112074 35460 112084
rect 35196 110572 35460 110582
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35196 110506 35460 110516
rect 35196 109004 35460 109014
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35196 108938 35460 108948
rect 35196 107436 35460 107446
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35196 107370 35460 107380
rect 35196 105868 35460 105878
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35196 105802 35460 105812
rect 35196 104300 35460 104310
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35196 104234 35460 104244
rect 35196 102732 35460 102742
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35196 102666 35460 102676
rect 35196 101164 35460 101174
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35196 101098 35460 101108
rect 35196 99596 35460 99606
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35196 99530 35460 99540
rect 35196 98028 35460 98038
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35196 97962 35460 97972
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 36652 66388 36708 114942
rect 37772 115556 37828 115566
rect 36652 66322 36708 66332
rect 36876 69972 36932 69982
rect 36876 65156 36932 69916
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 36876 65090 36932 65100
rect 35196 65034 35460 65044
rect 36316 64708 36372 64718
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 36316 57652 36372 64652
rect 37772 64036 37828 115500
rect 38668 115556 38724 115566
rect 38668 115462 38724 115500
rect 39788 102508 39844 116510
rect 41132 116340 41188 117070
rect 40796 116338 41188 116340
rect 40796 116286 41134 116338
rect 41186 116286 41188 116338
rect 40796 116284 41188 116286
rect 40796 115890 40852 116284
rect 41132 116274 41188 116284
rect 40796 115838 40798 115890
rect 40850 115838 40852 115890
rect 40796 115826 40852 115838
rect 41804 115892 41860 119200
rect 43148 116340 43204 119200
rect 43148 116274 43204 116284
rect 43484 116452 43540 116462
rect 42140 116004 42196 116014
rect 41916 115892 41972 115902
rect 41804 115890 41972 115892
rect 41804 115838 41918 115890
rect 41970 115838 41972 115890
rect 41804 115836 41972 115838
rect 41916 115826 41972 115836
rect 39452 102452 39844 102508
rect 41132 115556 41188 115566
rect 37884 99876 37940 99886
rect 37884 99316 37940 99820
rect 38556 99428 38612 99438
rect 38556 99334 38612 99372
rect 39452 99428 39508 102452
rect 38332 99316 38388 99326
rect 37884 99314 38388 99316
rect 37884 99262 37886 99314
rect 37938 99262 38334 99314
rect 38386 99262 38388 99314
rect 37884 99260 38388 99262
rect 37884 99250 37940 99260
rect 38332 99250 38388 99260
rect 39452 99314 39508 99372
rect 39452 99262 39454 99314
rect 39506 99262 39508 99314
rect 39452 99250 39508 99262
rect 39564 101780 39620 101790
rect 38892 99204 38948 99214
rect 38892 99110 38948 99148
rect 37772 63970 37828 63980
rect 36316 57586 36372 57596
rect 37772 60228 37828 60238
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 36204 56420 36260 56430
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 33964 53118 33966 53170
rect 34018 53118 34020 53170
rect 33964 53106 34020 53118
rect 33740 52946 33796 52958
rect 33740 52894 33742 52946
rect 33794 52894 33796 52946
rect 33740 52836 33796 52894
rect 34412 52836 34468 52846
rect 33740 52834 34468 52836
rect 33740 52782 34414 52834
rect 34466 52782 34468 52834
rect 33740 52780 34468 52782
rect 33516 52098 33572 52108
rect 34412 51156 34468 52780
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34412 51090 34468 51100
rect 34636 51156 34692 51166
rect 32732 47572 32788 47582
rect 32732 41188 32788 47516
rect 32732 41122 32788 41132
rect 32172 40404 32228 40414
rect 32172 4564 32228 40348
rect 34636 31220 34692 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 36092 40292 36148 40302
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34636 31154 34692 31164
rect 34412 31108 34468 31118
rect 32844 4564 32900 4574
rect 32172 4562 32900 4564
rect 32172 4510 32846 4562
rect 32898 4510 32900 4562
rect 32172 4508 32900 4510
rect 32172 4338 32228 4508
rect 32844 4498 32900 4508
rect 32172 4286 32174 4338
rect 32226 4286 32228 4338
rect 32172 4274 32228 4286
rect 31052 3614 31054 3666
rect 31106 3614 31108 3666
rect 26796 3602 26852 3612
rect 31052 3602 31108 3614
rect 31276 4226 31332 4238
rect 31276 4174 31278 4226
rect 31330 4174 31332 4226
rect 29372 3444 29428 3454
rect 29932 3444 29988 3454
rect 29372 3442 29988 3444
rect 29372 3390 29374 3442
rect 29426 3390 29934 3442
rect 29986 3390 29988 3442
rect 29372 3388 29988 3390
rect 29372 3378 29428 3388
rect 27692 3330 27748 3342
rect 27692 3278 27694 3330
rect 27746 3278 27748 3330
rect 27692 800 27748 3278
rect 28476 3332 28532 3342
rect 28476 3330 28868 3332
rect 28476 3278 28478 3330
rect 28530 3278 28868 3330
rect 28476 3276 28868 3278
rect 28476 3266 28532 3276
rect 24136 200 24360 728
rect 24444 700 24724 756
rect 24808 728 25060 800
rect 26152 728 26404 800
rect 27496 728 27748 800
rect 28812 800 28868 3276
rect 29484 800 29540 3388
rect 29932 3378 29988 3388
rect 31276 868 31332 4174
rect 34412 3780 34468 31052
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34524 21476 34580 21486
rect 34524 5236 34580 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34524 5170 34580 5180
rect 36092 5124 36148 40236
rect 36204 32452 36260 56364
rect 37548 41748 37604 41758
rect 37548 36596 37604 41692
rect 37772 40404 37828 60172
rect 39564 50372 39620 101724
rect 41132 67228 41188 115500
rect 42140 113428 42196 115948
rect 42140 113362 42196 113372
rect 41692 99204 41748 99214
rect 41132 67172 41300 67228
rect 41132 57090 41188 57102
rect 41132 57038 41134 57090
rect 41186 57038 41188 57090
rect 41132 56980 41188 57038
rect 40908 56978 41188 56980
rect 40908 56926 41134 56978
rect 41186 56926 41188 56978
rect 40908 56924 41188 56926
rect 40908 55522 40964 56924
rect 41132 56914 41188 56924
rect 40908 55470 40910 55522
rect 40962 55470 40964 55522
rect 40012 55412 40068 55422
rect 40012 55318 40068 55356
rect 40908 55412 40964 55470
rect 40796 55300 40852 55310
rect 40796 55206 40852 55244
rect 39676 55076 39732 55086
rect 39676 54982 39732 55020
rect 40684 55076 40740 55086
rect 40684 54982 40740 55020
rect 40796 54740 40852 54750
rect 40908 54740 40964 55356
rect 40796 54738 40964 54740
rect 40796 54686 40798 54738
rect 40850 54686 40964 54738
rect 40796 54684 40964 54686
rect 40796 54674 40852 54684
rect 40908 54628 40964 54684
rect 40908 54562 40964 54572
rect 40348 54404 40404 54414
rect 40348 54310 40404 54348
rect 39564 50306 39620 50316
rect 37772 40338 37828 40348
rect 39116 48804 39172 48814
rect 37548 36530 37604 36540
rect 36204 32386 36260 32396
rect 37772 33460 37828 33470
rect 37772 9268 37828 33404
rect 37772 9202 37828 9212
rect 36092 5058 36148 5068
rect 36540 4226 36596 4238
rect 36540 4174 36542 4226
rect 36594 4174 36596 4226
rect 36540 4116 36596 4174
rect 37660 4228 37716 4238
rect 37660 4226 37828 4228
rect 37660 4174 37662 4226
rect 37714 4174 37828 4226
rect 37660 4172 37828 4174
rect 37660 4162 37716 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34412 3714 34468 3724
rect 35532 3666 35588 3678
rect 35532 3614 35534 3666
rect 35586 3614 35588 3666
rect 33180 3330 33236 3342
rect 33180 3278 33182 3330
rect 33234 3278 33236 3330
rect 31052 812 31332 868
rect 32396 812 32564 868
rect 31052 800 31108 812
rect 32396 800 32452 812
rect 28812 728 29064 800
rect 29484 728 29736 800
rect 24808 200 25032 728
rect 26152 200 26376 728
rect 27496 200 27720 728
rect 28840 200 29064 728
rect 29512 200 29736 728
rect 30856 728 31108 800
rect 32200 728 32452 800
rect 32508 756 32564 812
rect 33180 756 33236 3278
rect 35532 800 35588 3614
rect 36316 3556 36372 3566
rect 36540 3556 36596 4060
rect 36316 3554 36596 3556
rect 36316 3502 36318 3554
rect 36370 3502 36596 3554
rect 36316 3500 36596 3502
rect 36316 3490 36372 3500
rect 37772 3444 37828 4172
rect 39116 3666 39172 48748
rect 41244 47796 41300 67172
rect 41468 57092 41524 57102
rect 41692 57092 41748 99148
rect 41468 57090 41748 57092
rect 41468 57038 41470 57090
rect 41522 57038 41748 57090
rect 41468 57036 41748 57038
rect 41468 57026 41524 57036
rect 41692 56866 41748 57036
rect 41692 56814 41694 56866
rect 41746 56814 41748 56866
rect 41692 56802 41748 56814
rect 42252 56754 42308 56766
rect 42252 56702 42254 56754
rect 42306 56702 42308 56754
rect 41692 55860 41748 55870
rect 41692 54738 41748 55804
rect 42252 55076 42308 56702
rect 42252 55010 42308 55020
rect 43372 55076 43428 55086
rect 41692 54686 41694 54738
rect 41746 54686 41748 54738
rect 41692 54674 41748 54686
rect 41580 54628 41636 54638
rect 41580 54534 41636 54572
rect 41804 54626 41860 54638
rect 41804 54574 41806 54626
rect 41858 54574 41860 54626
rect 41804 54404 41860 54574
rect 41804 54338 41860 54348
rect 42476 53844 42532 53854
rect 42476 53170 42532 53788
rect 42476 53118 42478 53170
rect 42530 53118 42532 53170
rect 42476 53106 42532 53118
rect 43372 53844 43428 55020
rect 43148 53058 43204 53070
rect 43148 53006 43150 53058
rect 43202 53006 43204 53058
rect 42028 52834 42084 52846
rect 42028 52782 42030 52834
rect 42082 52782 42084 52834
rect 42028 52052 42084 52782
rect 42028 51986 42084 51996
rect 43148 52052 43204 53006
rect 43372 53058 43428 53788
rect 43372 53006 43374 53058
rect 43426 53006 43428 53058
rect 43372 52994 43428 53006
rect 43260 52834 43316 52846
rect 43260 52782 43262 52834
rect 43314 52782 43316 52834
rect 43260 52052 43316 52782
rect 43372 52052 43428 52062
rect 43260 51996 43372 52052
rect 43148 51986 43204 51996
rect 43372 51986 43428 51996
rect 43484 48468 43540 116396
rect 43596 116226 43652 116238
rect 43596 116174 43598 116226
rect 43650 116174 43652 116226
rect 43596 116116 43652 116174
rect 43596 116050 43652 116060
rect 43596 115780 43652 115790
rect 43708 115780 43764 119200
rect 45052 116562 45108 119200
rect 45052 116510 45054 116562
rect 45106 116510 45108 116562
rect 44044 116340 44100 116350
rect 44044 116246 44100 116284
rect 43596 115778 43764 115780
rect 43596 115726 43598 115778
rect 43650 115726 43764 115778
rect 43596 115724 43764 115726
rect 45052 115780 45108 116510
rect 45388 115780 45444 115790
rect 45052 115778 45444 115780
rect 45052 115726 45390 115778
rect 45442 115726 45444 115778
rect 45052 115724 45444 115726
rect 43596 114996 43652 115724
rect 45388 115714 45444 115724
rect 46508 115780 46564 119200
rect 47628 119200 47880 119336
rect 48328 119200 48552 119800
rect 49672 119336 49896 119800
rect 49644 119200 49896 119336
rect 51016 119336 51240 119800
rect 51016 119200 51268 119336
rect 52360 119200 52584 119800
rect 53032 119336 53256 119800
rect 53032 119200 53284 119336
rect 54376 119200 54600 119800
rect 55720 119336 55944 119800
rect 56392 119336 56616 119800
rect 55692 119200 55944 119336
rect 56364 119200 56616 119336
rect 57736 119336 57960 119800
rect 59080 119336 59304 119800
rect 57736 119200 57988 119336
rect 59080 119200 59332 119336
rect 60424 119200 60648 119800
rect 61096 119200 61320 119800
rect 62440 119336 62664 119800
rect 63784 119336 64008 119800
rect 65128 119336 65352 119800
rect 62440 119200 62692 119336
rect 63784 119200 64036 119336
rect 65128 119200 65380 119336
rect 65800 119200 66024 119800
rect 67144 119336 67368 119800
rect 68488 119336 68712 119800
rect 67144 119200 67396 119336
rect 68488 119200 68740 119336
rect 69160 119200 69384 119800
rect 70504 119200 70728 119800
rect 71848 119336 72072 119800
rect 73192 119336 73416 119800
rect 71848 119200 72100 119336
rect 73192 119200 73444 119336
rect 73864 119200 74088 119800
rect 75208 119336 75432 119800
rect 76552 119336 76776 119800
rect 77896 119336 78120 119800
rect 78568 119336 78792 119800
rect 75208 119200 75460 119336
rect 76552 119200 76804 119336
rect 77896 119200 78148 119336
rect 78568 119200 78820 119336
rect 79912 119200 80136 119800
rect 81256 119336 81480 119800
rect 81928 119336 82152 119800
rect 81228 119200 81480 119336
rect 81900 119200 82152 119336
rect 83272 119336 83496 119800
rect 84616 119336 84840 119800
rect 85960 119336 86184 119800
rect 86632 119336 86856 119800
rect 87976 119336 88200 119800
rect 83272 119200 83524 119336
rect 84616 119200 84868 119336
rect 85960 119200 86212 119336
rect 86632 119200 86884 119336
rect 87976 119200 88228 119336
rect 89320 119200 89544 119800
rect 90664 119336 90888 119800
rect 90664 119200 90916 119336
rect 91336 119200 91560 119800
rect 92680 119200 92904 119800
rect 94024 119336 94248 119800
rect 94696 119336 94920 119800
rect 94024 119200 94276 119336
rect 94696 119200 94948 119336
rect 96040 119200 96264 119800
rect 97384 119336 97608 119800
rect 97384 119200 97636 119336
rect 98728 119200 98952 119800
rect 99400 119336 99624 119800
rect 99372 119200 99624 119336
rect 100744 119336 100968 119800
rect 100744 119200 100996 119336
rect 102088 119200 102312 119800
rect 102760 119200 102984 119800
rect 104104 119200 104328 119800
rect 105448 119200 105672 119800
rect 106792 119200 107016 119800
rect 107464 119200 107688 119800
rect 108808 119336 109032 119800
rect 108780 119200 109032 119336
rect 110152 119336 110376 119800
rect 110152 119200 110404 119336
rect 46956 116340 47012 116350
rect 46956 116246 47012 116284
rect 47628 116340 47684 119200
rect 47628 116274 47684 116284
rect 48076 116562 48132 116574
rect 48076 116510 48078 116562
rect 48130 116510 48132 116562
rect 48076 116228 48132 116510
rect 49532 116564 49588 116574
rect 49644 116564 49700 119200
rect 51212 117572 51268 119200
rect 51212 117516 51380 117572
rect 49532 116562 50148 116564
rect 49532 116510 49534 116562
rect 49586 116510 50148 116562
rect 49532 116508 50148 116510
rect 49532 116498 49588 116508
rect 48748 116340 48804 116350
rect 48748 116246 48804 116284
rect 50092 116338 50148 116508
rect 51212 116562 51268 116574
rect 51212 116510 51214 116562
rect 51266 116510 51268 116562
rect 51212 116452 51268 116510
rect 51212 116386 51268 116396
rect 50092 116286 50094 116338
rect 50146 116286 50148 116338
rect 50092 116274 50148 116286
rect 48076 116162 48132 116172
rect 48524 116116 48580 116126
rect 46508 115714 46564 115724
rect 47964 115780 48020 115790
rect 47292 115668 47348 115678
rect 46956 115666 47348 115668
rect 46956 115614 47294 115666
rect 47346 115614 47348 115666
rect 46956 115612 47348 115614
rect 43596 114930 43652 114940
rect 44492 115554 44548 115566
rect 44492 115502 44494 115554
rect 44546 115502 44548 115554
rect 44492 62188 44548 115502
rect 46508 115554 46564 115566
rect 46508 115502 46510 115554
rect 46562 115502 46564 115554
rect 45388 114996 45444 115006
rect 45388 114902 45444 114940
rect 46396 114996 46452 115006
rect 45276 105812 45332 105822
rect 44828 103234 44884 103246
rect 44828 103182 44830 103234
rect 44882 103182 44884 103234
rect 44828 103012 44884 103182
rect 44828 102946 44884 102956
rect 45164 103122 45220 103134
rect 45164 103070 45166 103122
rect 45218 103070 45220 103122
rect 45164 103012 45220 103070
rect 45164 102946 45220 102956
rect 44604 66500 44660 66510
rect 44604 65378 44660 66444
rect 44604 65326 44606 65378
rect 44658 65326 44660 65378
rect 44604 64820 44660 65326
rect 44716 64820 44772 64830
rect 44604 64818 44772 64820
rect 44604 64766 44718 64818
rect 44770 64766 44772 64818
rect 44604 64764 44772 64766
rect 44716 64596 44772 64764
rect 44716 64530 44772 64540
rect 44492 62132 44660 62188
rect 44492 58212 44548 58222
rect 44492 56308 44548 58156
rect 44604 57316 44660 62132
rect 45276 60116 45332 105756
rect 45612 103012 45668 103022
rect 45612 102918 45668 102956
rect 45948 103012 46004 103022
rect 45948 67228 46004 102956
rect 46396 68850 46452 114940
rect 46508 105812 46564 115502
rect 46956 114996 47012 115612
rect 47292 115602 47348 115612
rect 47964 115554 48020 115724
rect 47964 115502 47966 115554
rect 48018 115502 48020 115554
rect 47964 115490 48020 115502
rect 46956 114864 47012 114940
rect 46508 105746 46564 105756
rect 48300 93826 48356 93838
rect 48300 93774 48302 93826
rect 48354 93774 48356 93826
rect 48300 93604 48356 93774
rect 48300 93538 48356 93548
rect 46396 68798 46398 68850
rect 46450 68798 46452 68850
rect 46396 68786 46452 68798
rect 46060 68626 46116 68638
rect 46060 68574 46062 68626
rect 46114 68574 46116 68626
rect 46060 68516 46116 68574
rect 46060 68450 46116 68460
rect 46844 68516 46900 68526
rect 45724 67172 46004 67228
rect 45612 66274 45668 66286
rect 45612 66222 45614 66274
rect 45666 66222 45668 66274
rect 45612 64930 45668 66222
rect 45612 64878 45614 64930
rect 45666 64878 45668 64930
rect 45612 64866 45668 64878
rect 45612 63924 45668 63934
rect 45500 62354 45556 62366
rect 45500 62302 45502 62354
rect 45554 62302 45556 62354
rect 45500 61348 45556 62302
rect 45612 61570 45668 63868
rect 45724 63588 45780 67172
rect 46396 66724 46452 66734
rect 45836 66050 45892 66062
rect 45836 65998 45838 66050
rect 45890 65998 45892 66050
rect 45836 65604 45892 65998
rect 45836 65538 45892 65548
rect 45948 64708 46004 64718
rect 45948 64614 46004 64652
rect 45836 64036 45892 64046
rect 45836 63810 45892 63980
rect 45836 63758 45838 63810
rect 45890 63758 45892 63810
rect 45836 63746 45892 63758
rect 45724 62244 45780 63532
rect 45836 62468 45892 62478
rect 45836 62466 46340 62468
rect 45836 62414 45838 62466
rect 45890 62414 46340 62466
rect 45836 62412 46340 62414
rect 45836 62402 45892 62412
rect 45724 62188 46116 62244
rect 45612 61518 45614 61570
rect 45666 61518 45668 61570
rect 45612 61506 45668 61518
rect 45500 61292 45780 61348
rect 45724 61010 45780 61292
rect 45724 60958 45726 61010
rect 45778 60958 45780 61010
rect 45724 60946 45780 60958
rect 46060 60788 46116 62188
rect 46284 61682 46340 62412
rect 46396 62188 46452 66668
rect 46732 65604 46788 65614
rect 46732 65510 46788 65548
rect 46732 64932 46788 64942
rect 46732 64706 46788 64876
rect 46844 64820 46900 68460
rect 48412 67060 48468 67070
rect 48412 66966 48468 67004
rect 47964 66948 48020 66958
rect 47292 66388 47348 66398
rect 47292 66294 47348 66332
rect 47516 65492 47572 65502
rect 47516 65398 47572 65436
rect 47964 65490 48020 66892
rect 47964 65438 47966 65490
rect 48018 65438 48020 65490
rect 46844 64754 46900 64764
rect 47628 64932 47684 64942
rect 46732 64654 46734 64706
rect 46786 64654 46788 64706
rect 46732 64642 46788 64654
rect 47180 64708 47236 64718
rect 46508 64596 46564 64606
rect 46508 64502 46564 64540
rect 46844 64596 46900 64606
rect 46396 62132 46564 62188
rect 46284 61630 46286 61682
rect 46338 61630 46340 61682
rect 46284 61618 46340 61630
rect 46060 60656 46116 60732
rect 46508 60786 46564 62132
rect 46508 60734 46510 60786
rect 46562 60734 46564 60786
rect 45276 60050 45332 60060
rect 44604 57250 44660 57260
rect 46508 59778 46564 60734
rect 46620 60898 46676 60910
rect 46620 60846 46622 60898
rect 46674 60846 46676 60898
rect 46620 59892 46676 60846
rect 46620 59826 46676 59836
rect 46508 59726 46510 59778
rect 46562 59726 46564 59778
rect 45948 56868 46004 56878
rect 45948 56866 46452 56868
rect 45948 56814 45950 56866
rect 46002 56814 46452 56866
rect 45948 56812 46452 56814
rect 45948 56802 46004 56812
rect 44492 56242 44548 56252
rect 44940 56644 44996 56654
rect 44940 55970 44996 56588
rect 46172 56642 46228 56654
rect 46172 56590 46174 56642
rect 46226 56590 46228 56642
rect 46172 56196 46228 56590
rect 46172 56130 46228 56140
rect 44940 55918 44942 55970
rect 44994 55918 44996 55970
rect 44940 54740 44996 55918
rect 44940 54674 44996 54684
rect 45612 55972 45668 55982
rect 45388 53620 45444 53630
rect 45388 53526 45444 53564
rect 45052 51492 45108 51502
rect 45052 51398 45108 51436
rect 45388 51492 45444 51502
rect 45388 50708 45444 51436
rect 45500 51266 45556 51278
rect 45500 51214 45502 51266
rect 45554 51214 45556 51266
rect 45500 51156 45556 51214
rect 45500 51090 45556 51100
rect 45612 51154 45668 55916
rect 46396 55522 46452 56812
rect 46396 55470 46398 55522
rect 46450 55470 46452 55522
rect 46396 55458 46452 55470
rect 46508 55300 46564 59726
rect 46732 55300 46788 55310
rect 46396 55244 46564 55300
rect 46620 55298 46788 55300
rect 46620 55246 46734 55298
rect 46786 55246 46788 55298
rect 46620 55244 46788 55246
rect 45836 55074 45892 55086
rect 45836 55022 45838 55074
rect 45890 55022 45892 55074
rect 45724 54740 45780 54750
rect 45724 54646 45780 54684
rect 45724 54516 45780 54526
rect 45724 53170 45780 54460
rect 45836 54290 45892 55022
rect 46172 54628 46228 54638
rect 46172 54534 46228 54572
rect 46396 54404 46452 55244
rect 46508 54852 46564 54862
rect 46508 54738 46564 54796
rect 46508 54686 46510 54738
rect 46562 54686 46564 54738
rect 46508 54628 46564 54686
rect 46508 54562 46564 54572
rect 45836 54238 45838 54290
rect 45890 54238 45892 54290
rect 45836 54226 45892 54238
rect 46172 54348 46452 54404
rect 45948 53732 46004 53742
rect 45948 53638 46004 53676
rect 45724 53118 45726 53170
rect 45778 53118 45780 53170
rect 45724 53106 45780 53118
rect 46060 52276 46116 52286
rect 46060 52182 46116 52220
rect 45612 51102 45614 51154
rect 45666 51102 45668 51154
rect 45612 51090 45668 51102
rect 45836 51380 45892 51390
rect 45500 50708 45556 50718
rect 45388 50706 45556 50708
rect 45388 50654 45502 50706
rect 45554 50654 45556 50706
rect 45388 50652 45556 50654
rect 45500 50642 45556 50652
rect 45836 50596 45892 51324
rect 46060 51266 46116 51278
rect 46060 51214 46062 51266
rect 46114 51214 46116 51266
rect 46060 50932 46116 51214
rect 46060 50866 46116 50876
rect 45836 50034 45892 50540
rect 46172 50428 46228 54348
rect 46620 54290 46676 55244
rect 46732 55234 46788 55244
rect 46844 54516 46900 64540
rect 47180 64484 47236 64652
rect 47292 64484 47348 64494
rect 47180 64482 47348 64484
rect 47180 64430 47294 64482
rect 47346 64430 47348 64482
rect 47180 64428 47348 64430
rect 47068 60788 47124 60798
rect 47068 60114 47124 60732
rect 47068 60062 47070 60114
rect 47122 60062 47124 60114
rect 47068 60050 47124 60062
rect 46956 56642 47012 56654
rect 46956 56590 46958 56642
rect 47010 56590 47012 56642
rect 46956 56084 47012 56590
rect 47068 56196 47124 56206
rect 47068 56102 47124 56140
rect 46956 56018 47012 56028
rect 46620 54238 46622 54290
rect 46674 54238 46676 54290
rect 46396 53508 46452 53518
rect 45836 49982 45838 50034
rect 45890 49982 45892 50034
rect 45836 49970 45892 49982
rect 45948 50372 46228 50428
rect 46284 53506 46452 53508
rect 46284 53454 46398 53506
rect 46450 53454 46452 53506
rect 46284 53452 46452 53454
rect 45500 49812 45556 49822
rect 45500 49718 45556 49756
rect 45052 49700 45108 49710
rect 45276 49700 45332 49710
rect 45052 49698 45276 49700
rect 45052 49646 45054 49698
rect 45106 49646 45276 49698
rect 45052 49644 45276 49646
rect 45052 49634 45108 49644
rect 43484 48402 43540 48412
rect 45276 48466 45332 49644
rect 45724 49028 45780 49038
rect 45724 48804 45780 48972
rect 45724 48710 45780 48748
rect 45276 48414 45278 48466
rect 45330 48414 45332 48466
rect 45276 48402 45332 48414
rect 45724 48356 45780 48366
rect 45724 48132 45780 48300
rect 41244 47730 41300 47740
rect 45500 48130 45780 48132
rect 45500 48078 45726 48130
rect 45778 48078 45780 48130
rect 45500 48076 45780 48078
rect 45500 47572 45556 48076
rect 45724 48066 45780 48076
rect 45500 47478 45556 47516
rect 42924 46228 42980 46238
rect 42924 45332 42980 46172
rect 45612 46002 45668 46014
rect 45612 45950 45614 46002
rect 45666 45950 45668 46002
rect 42476 45330 42980 45332
rect 42476 45278 42926 45330
rect 42978 45278 42980 45330
rect 42476 45276 42980 45278
rect 42140 45220 42196 45230
rect 42140 45126 42196 45164
rect 42476 45218 42532 45276
rect 42924 45266 42980 45276
rect 43596 45556 43652 45566
rect 42476 45166 42478 45218
rect 42530 45166 42532 45218
rect 42476 45154 42532 45166
rect 41916 45108 41972 45118
rect 41132 43204 41188 43214
rect 39452 21364 39508 21374
rect 39452 20690 39508 21308
rect 39788 20916 39844 20926
rect 39788 20802 39844 20860
rect 40236 20916 40292 20926
rect 40236 20822 40292 20860
rect 41132 20916 41188 43148
rect 41916 42868 41972 45052
rect 41916 42802 41972 42812
rect 39788 20750 39790 20802
rect 39842 20750 39844 20802
rect 39788 20738 39844 20750
rect 39452 20638 39454 20690
rect 39506 20638 39508 20690
rect 39452 20626 39508 20638
rect 41132 20188 41188 20860
rect 43148 40628 43204 40638
rect 41132 20132 41636 20188
rect 41580 5236 41636 20132
rect 41580 5122 41636 5180
rect 41580 5070 41582 5122
rect 41634 5070 41636 5122
rect 41580 5058 41636 5070
rect 42028 5794 42084 5806
rect 42028 5742 42030 5794
rect 42082 5742 42084 5794
rect 40684 5012 40740 5022
rect 39116 3614 39118 3666
rect 39170 3614 39172 3666
rect 39116 3602 39172 3614
rect 40460 5010 40740 5012
rect 40460 4958 40686 5010
rect 40738 4958 40740 5010
rect 40460 4956 40740 4958
rect 37996 3444 38052 3454
rect 37772 3442 38052 3444
rect 37772 3390 37998 3442
rect 38050 3390 38052 3442
rect 37772 3388 38052 3390
rect 37212 3332 37268 3342
rect 37100 3330 37268 3332
rect 37100 3278 37214 3330
rect 37266 3278 37268 3330
rect 37100 3276 37268 3278
rect 37100 800 37156 3276
rect 37212 3266 37268 3276
rect 37772 800 37828 3388
rect 37996 3378 38052 3388
rect 40460 800 40516 4956
rect 40684 4946 40740 4956
rect 42028 4564 42084 5742
rect 42028 4498 42084 4508
rect 42364 5012 42420 5022
rect 42364 4564 42420 4956
rect 42364 4498 42420 4508
rect 42700 4898 42756 4910
rect 42700 4846 42702 4898
rect 42754 4846 42756 4898
rect 42700 4340 42756 4846
rect 43148 4676 43204 40572
rect 43596 6692 43652 45500
rect 45612 45108 45668 45950
rect 45612 45042 45668 45052
rect 44940 41860 44996 41870
rect 44940 31948 44996 41804
rect 45836 40292 45892 40302
rect 45836 40198 45892 40236
rect 45948 37044 46004 50372
rect 46284 49140 46340 53452
rect 46396 53442 46452 53452
rect 46620 52386 46676 54238
rect 46620 52334 46622 52386
rect 46674 52334 46676 52386
rect 46620 52322 46676 52334
rect 46732 54460 46900 54516
rect 46396 52162 46452 52174
rect 46396 52110 46398 52162
rect 46450 52110 46452 52162
rect 46396 51380 46452 52110
rect 46396 51314 46452 51324
rect 46508 51266 46564 51278
rect 46508 51214 46510 51266
rect 46562 51214 46564 51266
rect 46508 51154 46564 51214
rect 46508 51102 46510 51154
rect 46562 51102 46564 51154
rect 46508 51090 46564 51102
rect 46396 50484 46452 50494
rect 46396 50372 46452 50428
rect 46396 50034 46452 50316
rect 46396 49982 46398 50034
rect 46450 49982 46452 50034
rect 46396 49970 46452 49982
rect 46732 49810 46788 54460
rect 47068 54404 47124 54414
rect 46844 53956 46900 53966
rect 46844 53842 46900 53900
rect 46844 53790 46846 53842
rect 46898 53790 46900 53842
rect 46844 53778 46900 53790
rect 47068 53060 47124 54348
rect 47180 53284 47236 64428
rect 47292 64418 47348 64428
rect 47628 63138 47684 64876
rect 47964 64932 48020 65438
rect 47964 64866 48020 64876
rect 47852 64596 47908 64606
rect 47852 64502 47908 64540
rect 48188 64594 48244 64606
rect 48188 64542 48190 64594
rect 48242 64542 48244 64594
rect 47964 64482 48020 64494
rect 47964 64430 47966 64482
rect 48018 64430 48020 64482
rect 47964 64034 48020 64430
rect 48188 64484 48244 64542
rect 48188 64418 48244 64428
rect 48412 64594 48468 64606
rect 48412 64542 48414 64594
rect 48466 64542 48468 64594
rect 47964 63982 47966 64034
rect 48018 63982 48020 64034
rect 47964 63970 48020 63982
rect 48412 63812 48468 64542
rect 48412 63746 48468 63756
rect 47628 63086 47630 63138
rect 47682 63086 47684 63138
rect 47628 62188 47684 63086
rect 48188 63700 48244 63710
rect 48076 63026 48132 63038
rect 48076 62974 48078 63026
rect 48130 62974 48132 63026
rect 48076 62468 48132 62974
rect 47628 62132 47796 62188
rect 47740 60786 47796 62076
rect 47740 60734 47742 60786
rect 47794 60734 47796 60786
rect 47404 59892 47460 59902
rect 47404 59798 47460 59836
rect 47740 57540 47796 60734
rect 47964 60116 48020 60126
rect 47964 60022 48020 60060
rect 47852 57540 47908 57550
rect 47516 57538 47908 57540
rect 47516 57486 47854 57538
rect 47906 57486 47908 57538
rect 47516 57484 47908 57486
rect 47404 56868 47460 56878
rect 47404 56774 47460 56812
rect 47516 55298 47572 57484
rect 47852 57474 47908 57484
rect 47964 56642 48020 56654
rect 47964 56590 47966 56642
rect 48018 56590 48020 56642
rect 47852 56084 47908 56094
rect 47852 55990 47908 56028
rect 47964 55748 48020 56590
rect 47964 55682 48020 55692
rect 47516 55246 47518 55298
rect 47570 55246 47572 55298
rect 47516 55234 47572 55246
rect 47292 55186 47348 55198
rect 48076 55188 48132 62412
rect 48188 60674 48244 63644
rect 48300 62242 48356 62254
rect 48300 62190 48302 62242
rect 48354 62190 48356 62242
rect 48300 62132 48356 62190
rect 48300 62066 48356 62076
rect 48524 62020 48580 116060
rect 50556 116060 50820 116070
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50556 115994 50820 116004
rect 51324 115890 51380 117516
rect 52108 116676 52164 116686
rect 52108 116004 52164 116620
rect 53228 116564 53284 119200
rect 53228 116498 53284 116508
rect 54012 116564 54068 116574
rect 54012 116470 54068 116508
rect 53340 116450 53396 116462
rect 53340 116398 53342 116450
rect 53394 116398 53396 116450
rect 52780 116228 52836 116238
rect 53340 116228 53396 116398
rect 52108 115938 52164 115948
rect 52668 116226 53396 116228
rect 52668 116174 52782 116226
rect 52834 116174 53396 116226
rect 52668 116172 53396 116174
rect 51324 115838 51326 115890
rect 51378 115838 51380 115890
rect 51324 115826 51380 115838
rect 50556 114492 50820 114502
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50556 114426 50820 114436
rect 50556 112924 50820 112934
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50556 112858 50820 112868
rect 50556 111356 50820 111366
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50556 111290 50820 111300
rect 50556 109788 50820 109798
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50556 109722 50820 109732
rect 50556 108220 50820 108230
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50556 108154 50820 108164
rect 50556 106652 50820 106662
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50556 106586 50820 106596
rect 52444 105252 52500 105262
rect 50556 105084 50820 105094
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50556 105018 50820 105028
rect 50556 103516 50820 103526
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50556 103450 50820 103460
rect 50556 101948 50820 101958
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50556 101882 50820 101892
rect 50556 100380 50820 100390
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50556 100314 50820 100324
rect 50556 98812 50820 98822
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50556 98746 50820 98756
rect 50556 97244 50820 97254
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50556 97178 50820 97188
rect 50556 95676 50820 95686
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50556 95610 50820 95620
rect 50556 94108 50820 94118
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50556 94042 50820 94052
rect 48636 93714 48692 93726
rect 48636 93662 48638 93714
rect 48690 93662 48692 93714
rect 48636 93604 48692 93662
rect 48636 93538 48692 93548
rect 49420 93604 49476 93614
rect 49420 93510 49476 93548
rect 50556 92540 50820 92550
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50556 92474 50820 92484
rect 50556 90972 50820 90982
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50556 90906 50820 90916
rect 50556 89404 50820 89414
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50556 89338 50820 89348
rect 50556 87836 50820 87846
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50556 87770 50820 87780
rect 50556 86268 50820 86278
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50556 86202 50820 86212
rect 50556 84700 50820 84710
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50556 84634 50820 84644
rect 50556 83132 50820 83142
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50556 83066 50820 83076
rect 50556 81564 50820 81574
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50556 81498 50820 81508
rect 50556 79996 50820 80006
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50556 79930 50820 79940
rect 50556 78428 50820 78438
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50556 78362 50820 78372
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 49308 67844 49364 67854
rect 49308 67842 49812 67844
rect 49308 67790 49310 67842
rect 49362 67790 49812 67842
rect 49308 67788 49812 67790
rect 49308 67778 49364 67788
rect 49644 67618 49700 67630
rect 49644 67566 49646 67618
rect 49698 67566 49700 67618
rect 49644 67228 49700 67566
rect 48636 67170 48692 67182
rect 48636 67118 48638 67170
rect 48690 67118 48692 67170
rect 48636 66388 48692 67118
rect 49532 67172 49700 67228
rect 49532 66500 49588 67116
rect 49644 67060 49700 67070
rect 49644 66966 49700 67004
rect 49532 66434 49588 66444
rect 49756 66836 49812 67788
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50540 67172 50596 67182
rect 50540 67078 50596 67116
rect 50764 67058 50820 67070
rect 50764 67006 50766 67058
rect 50818 67006 50820 67058
rect 50764 66948 50820 67006
rect 51996 67060 52052 67070
rect 49980 66836 50036 66846
rect 49756 66834 50036 66836
rect 49756 66782 49982 66834
rect 50034 66782 50036 66834
rect 49756 66780 50036 66782
rect 48636 66322 48692 66332
rect 49420 66388 49476 66398
rect 49420 66294 49476 66332
rect 48636 65492 48692 65502
rect 48636 63924 48692 65436
rect 49532 65492 49588 65502
rect 49532 65398 49588 65436
rect 48748 65378 48804 65390
rect 48748 65326 48750 65378
rect 48802 65326 48804 65378
rect 48748 65268 48804 65326
rect 48748 64596 48804 65212
rect 48748 64530 48804 64540
rect 49196 64482 49252 64494
rect 49196 64430 49198 64482
rect 49250 64430 49252 64482
rect 48692 63868 48916 63924
rect 48636 63792 48692 63868
rect 48636 63252 48692 63262
rect 48636 63158 48692 63196
rect 48524 61954 48580 61964
rect 48860 62244 48916 63868
rect 49196 62468 49252 64430
rect 49644 64482 49700 64494
rect 49644 64430 49646 64482
rect 49698 64430 49700 64482
rect 49644 64036 49700 64430
rect 49644 63942 49700 63980
rect 49532 63812 49588 63822
rect 49532 63718 49588 63756
rect 49196 62402 49252 62412
rect 49532 62468 49588 62478
rect 49532 62374 49588 62412
rect 49756 62244 49812 66780
rect 49980 66770 50036 66780
rect 50764 66724 50820 66892
rect 50764 66658 50820 66668
rect 51324 66946 51380 66958
rect 51324 66894 51326 66946
rect 51378 66894 51380 66946
rect 51324 66724 51380 66894
rect 51324 66658 51380 66668
rect 50204 66332 50708 66388
rect 50204 66274 50260 66332
rect 50204 66222 50206 66274
rect 50258 66222 50260 66274
rect 50204 66210 50260 66222
rect 50652 66052 50708 66332
rect 50652 65986 50708 65996
rect 51884 66164 51940 66174
rect 51884 66050 51940 66108
rect 51884 65998 51886 66050
rect 51938 65998 51940 66050
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 49980 65492 50036 65502
rect 49980 65398 50036 65436
rect 50204 64482 50260 64494
rect 50204 64430 50206 64482
rect 50258 64430 50260 64482
rect 49868 63698 49924 63710
rect 49868 63646 49870 63698
rect 49922 63646 49924 63698
rect 49868 62916 49924 63646
rect 50204 63700 50260 64430
rect 50652 64484 50708 64522
rect 50652 64418 50708 64428
rect 51436 64484 51492 64494
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50764 63924 50820 63934
rect 51212 63924 51268 63934
rect 50764 63922 51268 63924
rect 50764 63870 50766 63922
rect 50818 63870 51214 63922
rect 51266 63870 51268 63922
rect 50764 63868 51268 63870
rect 50428 63812 50484 63822
rect 50428 63718 50484 63756
rect 50540 63810 50596 63822
rect 50540 63758 50542 63810
rect 50594 63758 50596 63810
rect 50204 63634 50260 63644
rect 49868 62468 49924 62860
rect 50316 63028 50372 63038
rect 50540 63028 50596 63758
rect 50764 63252 50820 63868
rect 51212 63858 51268 63868
rect 50764 63186 50820 63196
rect 50316 62578 50372 62972
rect 50316 62526 50318 62578
rect 50370 62526 50372 62578
rect 50316 62514 50372 62526
rect 50428 62972 50596 63028
rect 50764 63028 50820 63038
rect 50428 62580 50484 62972
rect 50764 62934 50820 62972
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 51324 62580 51380 62590
rect 50428 62524 50596 62580
rect 49868 62402 49924 62412
rect 50092 62468 50148 62478
rect 50092 62374 50148 62412
rect 48412 61684 48468 61694
rect 48860 61684 48916 62188
rect 49420 62188 49812 62244
rect 50428 62354 50484 62366
rect 50428 62302 50430 62354
rect 50482 62302 50484 62354
rect 48412 61682 48580 61684
rect 48412 61630 48414 61682
rect 48466 61630 48580 61682
rect 48412 61628 48580 61630
rect 48412 61618 48468 61628
rect 48188 60622 48190 60674
rect 48242 60622 48244 60674
rect 48188 55748 48244 60622
rect 48524 59892 48580 61628
rect 48748 61682 48916 61684
rect 48748 61630 48862 61682
rect 48914 61630 48916 61682
rect 48748 61628 48916 61630
rect 48748 60228 48804 61628
rect 48860 61618 48916 61628
rect 49308 62132 49364 62142
rect 49308 61682 49364 62076
rect 49308 61630 49310 61682
rect 49362 61630 49364 61682
rect 49308 61618 49364 61630
rect 49420 60228 49476 62188
rect 50428 62132 50484 62302
rect 50540 62354 50596 62524
rect 50540 62302 50542 62354
rect 50594 62302 50596 62354
rect 50540 62290 50596 62302
rect 51100 62354 51156 62366
rect 51100 62302 51102 62354
rect 51154 62302 51156 62354
rect 50428 62066 50484 62076
rect 51100 62132 51156 62302
rect 50428 61684 50484 61694
rect 50204 60788 50260 60798
rect 50204 60694 50260 60732
rect 49532 60676 49588 60686
rect 50316 60676 50372 60686
rect 49532 60674 49812 60676
rect 49532 60622 49534 60674
rect 49586 60622 49812 60674
rect 49532 60620 49812 60622
rect 49532 60610 49588 60620
rect 48524 59826 48580 59836
rect 48636 60172 48804 60228
rect 49308 60172 49476 60228
rect 48300 59778 48356 59790
rect 48300 59726 48302 59778
rect 48354 59726 48356 59778
rect 48300 59668 48356 59726
rect 48300 59602 48356 59612
rect 48412 58436 48468 58446
rect 48636 58436 48692 60172
rect 49196 60116 49252 60126
rect 49196 60022 49252 60060
rect 48748 60004 48804 60014
rect 48748 59910 48804 59948
rect 48972 59668 49028 59678
rect 48748 59220 48804 59230
rect 48748 59126 48804 59164
rect 48412 58434 48692 58436
rect 48412 58382 48414 58434
rect 48466 58382 48692 58434
rect 48412 58380 48692 58382
rect 48412 58370 48468 58380
rect 48412 57538 48468 57550
rect 48412 57486 48414 57538
rect 48466 57486 48468 57538
rect 48412 56420 48468 57486
rect 48412 56354 48468 56364
rect 48524 56866 48580 58380
rect 48524 56814 48526 56866
rect 48578 56814 48580 56866
rect 48524 56084 48580 56814
rect 48748 57540 48804 57550
rect 48524 56018 48580 56028
rect 48636 56196 48692 56206
rect 48300 55972 48356 55982
rect 48300 55878 48356 55916
rect 48188 55692 48580 55748
rect 47292 55134 47294 55186
rect 47346 55134 47348 55186
rect 47292 54740 47348 55134
rect 47292 54674 47348 54684
rect 47740 55132 48132 55188
rect 48300 55524 48356 55534
rect 47404 54516 47460 54526
rect 47404 53732 47460 54460
rect 47404 53666 47460 53676
rect 47292 53508 47348 53518
rect 47292 53414 47348 53452
rect 47628 53506 47684 53518
rect 47628 53454 47630 53506
rect 47682 53454 47684 53506
rect 47628 53396 47684 53454
rect 47180 53218 47236 53228
rect 47404 53340 47628 53396
rect 47068 53004 47348 53060
rect 47068 52500 47124 52510
rect 46956 51940 47012 51950
rect 46732 49758 46734 49810
rect 46786 49758 46788 49810
rect 46732 49700 46788 49758
rect 46508 49140 46564 49150
rect 46284 49084 46508 49140
rect 46508 49046 46564 49084
rect 46060 48916 46116 48926
rect 46060 48822 46116 48860
rect 46732 48354 46788 49644
rect 46844 51938 47012 51940
rect 46844 51886 46958 51938
rect 47010 51886 47012 51938
rect 46844 51884 47012 51886
rect 46844 50260 46900 51884
rect 46956 51874 47012 51884
rect 46956 51266 47012 51278
rect 46956 51214 46958 51266
rect 47010 51214 47012 51266
rect 46956 51156 47012 51214
rect 46956 51090 47012 51100
rect 47068 50428 47124 52444
rect 46844 49140 46900 50204
rect 46956 50372 47124 50428
rect 47292 52274 47348 53004
rect 47292 52222 47294 52274
rect 47346 52222 47348 52274
rect 46956 49812 47012 50372
rect 47068 50148 47124 50158
rect 47068 50034 47124 50092
rect 47068 49982 47070 50034
rect 47122 49982 47124 50034
rect 47068 49970 47124 49982
rect 47068 49812 47124 49822
rect 46956 49756 47068 49812
rect 47068 49718 47124 49756
rect 46956 49140 47012 49150
rect 46844 49138 47012 49140
rect 46844 49086 46958 49138
rect 47010 49086 47012 49138
rect 46844 49084 47012 49086
rect 46956 49074 47012 49084
rect 46732 48302 46734 48354
rect 46786 48302 46788 48354
rect 46284 48132 46340 48142
rect 46284 48038 46340 48076
rect 46732 46900 46788 48302
rect 47068 48804 47124 48814
rect 47292 48804 47348 52222
rect 47404 50708 47460 53340
rect 47628 53330 47684 53340
rect 47740 52836 47796 55132
rect 48188 55076 48244 55114
rect 48188 55010 48244 55020
rect 47852 54964 47908 54974
rect 47852 54738 47908 54908
rect 47852 54686 47854 54738
rect 47906 54686 47908 54738
rect 47852 54674 47908 54686
rect 48188 54852 48244 54862
rect 47964 54404 48020 54414
rect 47964 53620 48020 54348
rect 48188 53844 48244 54796
rect 48188 53778 48244 53788
rect 48188 53620 48244 53630
rect 47964 53618 48244 53620
rect 47964 53566 48190 53618
rect 48242 53566 48244 53618
rect 47964 53564 48244 53566
rect 48188 53554 48244 53564
rect 48076 53284 48132 53294
rect 47740 52780 47908 52836
rect 47740 52612 47796 52622
rect 47740 52274 47796 52556
rect 47740 52222 47742 52274
rect 47794 52222 47796 52274
rect 47740 52164 47796 52222
rect 47740 52098 47796 52108
rect 47852 52276 47908 52780
rect 47964 52834 48020 52846
rect 47964 52782 47966 52834
rect 48018 52782 48020 52834
rect 47964 52388 48020 52782
rect 47964 52322 48020 52332
rect 48076 52724 48132 53228
rect 47516 51492 47572 51502
rect 47516 51398 47572 51436
rect 47740 51492 47796 51502
rect 47852 51492 47908 52220
rect 48076 52164 48132 52668
rect 48188 52386 48244 52398
rect 48188 52334 48190 52386
rect 48242 52334 48244 52386
rect 48188 52274 48244 52334
rect 48188 52222 48190 52274
rect 48242 52222 48244 52274
rect 48188 52210 48244 52222
rect 48076 52098 48132 52108
rect 48300 51492 48356 55468
rect 48412 54402 48468 54414
rect 48412 54350 48414 54402
rect 48466 54350 48468 54402
rect 48412 54180 48468 54350
rect 48412 54114 48468 54124
rect 48412 53844 48468 53854
rect 48412 53730 48468 53788
rect 48412 53678 48414 53730
rect 48466 53678 48468 53730
rect 48412 53666 48468 53678
rect 48412 52500 48468 52510
rect 48412 52276 48468 52444
rect 48412 51602 48468 52220
rect 48412 51550 48414 51602
rect 48466 51550 48468 51602
rect 48412 51538 48468 51550
rect 47740 51490 47908 51492
rect 47740 51438 47742 51490
rect 47794 51438 47908 51490
rect 47740 51436 47908 51438
rect 48188 51436 48356 51492
rect 47740 51426 47796 51436
rect 47628 51266 47684 51278
rect 47628 51214 47630 51266
rect 47682 51214 47684 51266
rect 47628 50820 47684 51214
rect 48076 51268 48132 51278
rect 47628 50764 47908 50820
rect 47404 50652 47796 50708
rect 47628 50482 47684 50494
rect 47628 50430 47630 50482
rect 47682 50430 47684 50482
rect 47628 50428 47684 50430
rect 47516 50372 47684 50428
rect 47404 50316 47572 50372
rect 47404 50148 47460 50316
rect 47404 50082 47460 50092
rect 47740 50036 47796 50652
rect 47516 49980 47796 50036
rect 47404 49924 47460 49934
rect 47404 49830 47460 49868
rect 47404 48804 47460 48814
rect 47292 48802 47460 48804
rect 47292 48750 47406 48802
rect 47458 48750 47460 48802
rect 47292 48748 47460 48750
rect 47068 48354 47124 48748
rect 47404 48692 47460 48748
rect 47404 48626 47460 48636
rect 47516 48468 47572 49980
rect 47852 49924 47908 50764
rect 47964 50372 48020 50382
rect 47964 50034 48020 50316
rect 47964 49982 47966 50034
rect 48018 49982 48020 50034
rect 47964 49970 48020 49982
rect 47852 49858 47908 49868
rect 47852 49140 47908 49150
rect 47852 49046 47908 49084
rect 47068 48302 47070 48354
rect 47122 48302 47124 48354
rect 47068 48290 47124 48302
rect 47180 48412 47572 48468
rect 46844 48130 46900 48142
rect 46844 48078 46846 48130
rect 46898 48078 46900 48130
rect 46844 47572 46900 48078
rect 46844 47506 46900 47516
rect 46844 46900 46900 46910
rect 46732 46844 46844 46900
rect 46844 46768 46900 46844
rect 46956 45108 47012 45118
rect 46956 45014 47012 45052
rect 47068 44100 47124 44110
rect 45948 36978 46004 36988
rect 46620 37044 46676 37054
rect 45836 34916 45892 34926
rect 45836 34914 46004 34916
rect 45836 34862 45838 34914
rect 45890 34862 46004 34914
rect 45836 34860 46004 34862
rect 45836 34850 45892 34860
rect 45052 34020 45108 34030
rect 45108 33964 45332 34020
rect 45052 33926 45108 33964
rect 45276 33460 45332 33964
rect 45948 33572 46004 34860
rect 46060 34690 46116 34702
rect 46060 34638 46062 34690
rect 46114 34638 46116 34690
rect 46060 34244 46116 34638
rect 46060 34178 46116 34188
rect 46060 33572 46116 33582
rect 45948 33570 46116 33572
rect 45948 33518 46062 33570
rect 46114 33518 46116 33570
rect 45948 33516 46116 33518
rect 46060 33506 46116 33516
rect 45388 33460 45444 33470
rect 45276 33458 45444 33460
rect 45276 33406 45390 33458
rect 45442 33406 45444 33458
rect 45276 33404 45444 33406
rect 45388 33236 45444 33404
rect 46396 33460 46452 33470
rect 46396 33366 46452 33404
rect 45388 33170 45444 33180
rect 46620 33348 46676 36988
rect 46620 33234 46676 33292
rect 46620 33182 46622 33234
rect 46674 33182 46676 33234
rect 46620 33170 46676 33182
rect 46956 33236 47012 33246
rect 46956 33142 47012 33180
rect 47068 31948 47124 44044
rect 47180 38668 47236 48412
rect 47964 48356 48020 48366
rect 47964 48262 48020 48300
rect 47292 48242 47348 48254
rect 47292 48190 47294 48242
rect 47346 48190 47348 48242
rect 47292 48132 47348 48190
rect 47852 48132 47908 48142
rect 47292 48130 47908 48132
rect 47292 48078 47854 48130
rect 47906 48078 47908 48130
rect 47292 48076 47908 48078
rect 47852 48066 47908 48076
rect 48076 48020 48132 51212
rect 48188 50428 48244 51436
rect 48300 51268 48356 51278
rect 48300 51174 48356 51212
rect 48300 50596 48356 50634
rect 48300 50530 48356 50540
rect 48524 50428 48580 55692
rect 48636 55524 48692 56140
rect 48636 55458 48692 55468
rect 48636 55076 48692 55086
rect 48748 55076 48804 57484
rect 48860 56084 48916 56094
rect 48860 55990 48916 56028
rect 48972 55300 49028 59612
rect 49308 59332 49364 60172
rect 49644 60114 49700 60126
rect 49644 60062 49646 60114
rect 49698 60062 49700 60114
rect 49308 59220 49364 59276
rect 49196 59164 49364 59220
rect 49420 60004 49476 60014
rect 49084 58548 49140 58558
rect 49084 58454 49140 58492
rect 49196 56980 49252 59164
rect 48972 55234 49028 55244
rect 49084 56924 49252 56980
rect 48636 55074 48804 55076
rect 48636 55022 48638 55074
rect 48690 55022 48804 55074
rect 48636 55020 48804 55022
rect 48636 55010 48692 55020
rect 48636 54516 48692 54526
rect 48748 54516 48804 55020
rect 49084 54852 49140 56924
rect 49196 56754 49252 56766
rect 49196 56702 49198 56754
rect 49250 56702 49252 56754
rect 49196 55524 49252 56702
rect 49196 55458 49252 55468
rect 49196 55300 49252 55310
rect 49196 55206 49252 55244
rect 49084 54786 49140 54796
rect 49308 54964 49364 54974
rect 48860 54740 48916 54750
rect 48860 54646 48916 54684
rect 48748 54460 48916 54516
rect 48636 53618 48692 54460
rect 48748 53844 48804 53854
rect 48748 53750 48804 53788
rect 48636 53566 48638 53618
rect 48690 53566 48692 53618
rect 48636 53554 48692 53566
rect 48860 53508 48916 54460
rect 49196 53620 49252 53630
rect 49196 53526 49252 53564
rect 48860 53442 48916 53452
rect 49084 53396 49140 53406
rect 48748 52946 48804 52958
rect 48748 52894 48750 52946
rect 48802 52894 48804 52946
rect 48636 52500 48692 52510
rect 48636 52386 48692 52444
rect 48636 52334 48638 52386
rect 48690 52334 48692 52386
rect 48636 52322 48692 52334
rect 48636 52164 48692 52174
rect 48636 52070 48692 52108
rect 48748 51380 48804 52894
rect 49084 51940 49140 53340
rect 49196 52388 49252 52398
rect 49196 52294 49252 52332
rect 49084 51884 49252 51940
rect 48748 50596 48804 51324
rect 49084 51492 49140 51502
rect 48748 50530 48804 50540
rect 48972 51044 49028 51054
rect 48188 50372 48356 50428
rect 48524 50372 48692 50428
rect 48076 47954 48132 47964
rect 48188 48132 48244 48142
rect 48188 48018 48244 48076
rect 48188 47966 48190 48018
rect 48242 47966 48244 48018
rect 47628 47572 47684 47582
rect 47628 47478 47684 47516
rect 47292 46900 47348 46910
rect 47292 46786 47348 46844
rect 47292 46734 47294 46786
rect 47346 46734 47348 46786
rect 47292 46722 47348 46734
rect 47516 46898 47572 46910
rect 47516 46846 47518 46898
rect 47570 46846 47572 46898
rect 47516 46004 47572 46846
rect 47628 46676 47684 46686
rect 47628 46582 47684 46620
rect 47852 46674 47908 46686
rect 47852 46622 47854 46674
rect 47906 46622 47908 46674
rect 47740 46004 47796 46014
rect 47516 46002 47796 46004
rect 47516 45950 47742 46002
rect 47794 45950 47796 46002
rect 47516 45948 47796 45950
rect 47740 45938 47796 45948
rect 47740 45332 47796 45342
rect 47852 45332 47908 46622
rect 47740 45330 47908 45332
rect 47740 45278 47742 45330
rect 47794 45278 47908 45330
rect 47740 45276 47908 45278
rect 47740 45266 47796 45276
rect 47516 45108 47572 45118
rect 47516 45014 47572 45052
rect 47852 44884 47908 44894
rect 48188 44884 48244 47966
rect 47852 44882 48244 44884
rect 47852 44830 47854 44882
rect 47906 44830 48244 44882
rect 47852 44828 48244 44830
rect 47852 44100 47908 44828
rect 48300 44548 48356 50372
rect 48524 50036 48580 50046
rect 48412 49700 48468 49710
rect 48412 49606 48468 49644
rect 48412 49140 48468 49150
rect 48524 49140 48580 49980
rect 48412 49138 48580 49140
rect 48412 49086 48414 49138
rect 48466 49086 48580 49138
rect 48412 49084 48580 49086
rect 48412 49074 48468 49084
rect 48636 48132 48692 50372
rect 48748 50036 48804 50046
rect 48748 49942 48804 49980
rect 48860 49924 48916 49934
rect 48860 49138 48916 49868
rect 48860 49086 48862 49138
rect 48914 49086 48916 49138
rect 48860 49074 48916 49086
rect 48860 48468 48916 48478
rect 48972 48468 49028 50988
rect 48860 48466 49028 48468
rect 48860 48414 48862 48466
rect 48914 48414 49028 48466
rect 48860 48412 49028 48414
rect 49084 50932 49140 51436
rect 48860 48402 48916 48412
rect 48636 48066 48692 48076
rect 49084 47796 49140 50876
rect 49196 50706 49252 51884
rect 49196 50654 49198 50706
rect 49250 50654 49252 50706
rect 49196 50642 49252 50654
rect 49308 51938 49364 54908
rect 49308 51886 49310 51938
rect 49362 51886 49364 51938
rect 49308 50260 49364 51886
rect 49196 49700 49252 49710
rect 49196 48468 49252 49644
rect 49308 49364 49364 50204
rect 49308 49298 49364 49308
rect 49420 53730 49476 59948
rect 49532 59778 49588 59790
rect 49532 59726 49534 59778
rect 49586 59726 49588 59778
rect 49532 59330 49588 59726
rect 49644 59668 49700 60062
rect 49756 60002 49812 60620
rect 50316 60228 50372 60620
rect 49756 59950 49758 60002
rect 49810 59950 49812 60002
rect 49756 59938 49812 59950
rect 50092 60172 50372 60228
rect 49644 59602 49700 59612
rect 49532 59278 49534 59330
rect 49586 59278 49588 59330
rect 49532 59266 49588 59278
rect 49756 59330 49812 59342
rect 49756 59278 49758 59330
rect 49810 59278 49812 59330
rect 49756 59220 49812 59278
rect 49644 59106 49700 59118
rect 49644 59054 49646 59106
rect 49698 59054 49700 59106
rect 49644 58548 49700 59054
rect 49644 58482 49700 58492
rect 49532 57764 49588 57774
rect 49532 57670 49588 57708
rect 49644 56420 49700 56430
rect 49644 56194 49700 56364
rect 49644 56142 49646 56194
rect 49698 56142 49700 56194
rect 49644 56130 49700 56142
rect 49644 55524 49700 55562
rect 49644 55458 49700 55468
rect 49756 55074 49812 59164
rect 49868 57650 49924 57662
rect 49868 57598 49870 57650
rect 49922 57598 49924 57650
rect 49868 57540 49924 57598
rect 49868 57474 49924 57484
rect 50092 56532 50148 60172
rect 50204 60002 50260 60014
rect 50204 59950 50206 60002
rect 50258 59950 50260 60002
rect 50204 59892 50260 59950
rect 50316 60004 50372 60014
rect 50316 59910 50372 59948
rect 50428 60002 50484 61628
rect 50876 61346 50932 61358
rect 50876 61294 50878 61346
rect 50930 61294 50932 61346
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50428 59950 50430 60002
rect 50482 59950 50484 60002
rect 50428 59938 50484 59950
rect 50204 59826 50260 59836
rect 50876 59892 50932 61294
rect 51100 61124 51156 62076
rect 51324 62244 51380 62524
rect 51212 61684 51268 61694
rect 51212 61590 51268 61628
rect 51100 61058 51156 61068
rect 50876 59826 50932 59836
rect 50988 60788 51044 60798
rect 50988 60674 51044 60732
rect 50988 60622 50990 60674
rect 51042 60622 51044 60674
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50988 59556 51044 60622
rect 51212 60228 51268 60238
rect 50988 59490 51044 59500
rect 51100 60226 51268 60228
rect 51100 60174 51214 60226
rect 51266 60174 51268 60226
rect 51100 60172 51268 60174
rect 50764 59108 50820 59118
rect 51100 59108 51156 60172
rect 51212 60162 51268 60172
rect 51324 59780 51380 62188
rect 50764 59106 51156 59108
rect 50764 59054 50766 59106
rect 50818 59054 51156 59106
rect 50764 59052 51156 59054
rect 51212 59778 51380 59780
rect 51212 59726 51326 59778
rect 51378 59726 51380 59778
rect 51212 59724 51380 59726
rect 50764 59042 50820 59052
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50540 57540 50596 57550
rect 50540 57446 50596 57484
rect 50428 56868 50484 56878
rect 50092 56476 50372 56532
rect 50092 56308 50148 56318
rect 49980 56306 50148 56308
rect 49980 56254 50094 56306
rect 50146 56254 50148 56306
rect 49980 56252 50148 56254
rect 49868 55970 49924 55982
rect 49868 55918 49870 55970
rect 49922 55918 49924 55970
rect 49868 55748 49924 55918
rect 49868 55682 49924 55692
rect 49980 55522 50036 56252
rect 50092 56242 50148 56252
rect 50204 56084 50260 56094
rect 50204 55990 50260 56028
rect 49980 55470 49982 55522
rect 50034 55470 50036 55522
rect 49980 55458 50036 55470
rect 50092 55858 50148 55870
rect 50092 55806 50094 55858
rect 50146 55806 50148 55858
rect 50092 55524 50148 55806
rect 50316 55636 50372 56476
rect 50428 56308 50484 56812
rect 50876 56644 50932 59052
rect 50988 57540 51044 57550
rect 50988 57446 51044 57484
rect 51212 57540 51268 59724
rect 51324 59714 51380 59724
rect 51324 59556 51380 59566
rect 51324 58210 51380 59500
rect 51324 58158 51326 58210
rect 51378 58158 51380 58210
rect 51324 58100 51380 58158
rect 51324 58034 51380 58044
rect 51436 57764 51492 64428
rect 51772 63364 51828 63374
rect 51548 63362 51828 63364
rect 51548 63310 51774 63362
rect 51826 63310 51828 63362
rect 51548 63308 51828 63310
rect 51548 63138 51604 63308
rect 51772 63298 51828 63308
rect 51548 63086 51550 63138
rect 51602 63086 51604 63138
rect 51548 63074 51604 63086
rect 51548 60676 51604 60686
rect 51548 60582 51604 60620
rect 51884 60226 51940 65998
rect 51996 66052 52052 67004
rect 52332 66164 52388 66174
rect 52332 66070 52388 66108
rect 51996 63362 52052 65996
rect 51996 63310 51998 63362
rect 52050 63310 52052 63362
rect 51996 63250 52052 63310
rect 51996 63198 51998 63250
rect 52050 63198 52052 63250
rect 51996 63186 52052 63198
rect 52444 61684 52500 105196
rect 52668 90748 52724 116172
rect 52780 116162 52836 116172
rect 53116 116004 53172 116014
rect 52668 90692 52836 90748
rect 52668 67060 52724 67070
rect 52668 66966 52724 67004
rect 52668 66164 52724 66174
rect 52780 66164 52836 90692
rect 52668 66162 52836 66164
rect 52668 66110 52670 66162
rect 52722 66110 52836 66162
rect 52668 66108 52836 66110
rect 52668 66098 52724 66108
rect 52892 62356 52948 62366
rect 52892 62262 52948 62300
rect 52444 61618 52500 61628
rect 52220 61348 52276 61358
rect 52220 61254 52276 61292
rect 52668 61346 52724 61358
rect 52668 61294 52670 61346
rect 52722 61294 52724 61346
rect 52668 61236 52724 61294
rect 52668 61170 52724 61180
rect 52668 61012 52724 61022
rect 52668 60918 52724 60956
rect 51884 60174 51886 60226
rect 51938 60174 51940 60226
rect 51884 60162 51940 60174
rect 52220 60674 52276 60686
rect 52220 60622 52222 60674
rect 52274 60622 52276 60674
rect 51884 60004 51940 60014
rect 51884 59910 51940 59948
rect 51212 57474 51268 57484
rect 51324 57708 51492 57764
rect 51772 59892 51828 59902
rect 50876 56578 50932 56588
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50428 56252 50596 56308
rect 50540 56082 50596 56252
rect 51100 56196 51156 56206
rect 51100 56102 51156 56140
rect 50540 56030 50542 56082
rect 50594 56030 50596 56082
rect 50540 56018 50596 56030
rect 50652 56084 50708 56094
rect 50540 55860 50596 55870
rect 50652 55860 50708 56028
rect 50764 55860 50820 55870
rect 50652 55858 50820 55860
rect 50652 55806 50766 55858
rect 50818 55806 50820 55858
rect 50652 55804 50820 55806
rect 50540 55636 50596 55804
rect 50764 55794 50820 55804
rect 50652 55636 50708 55646
rect 50540 55580 50652 55636
rect 50316 55570 50372 55580
rect 50652 55570 50708 55580
rect 50092 55458 50148 55468
rect 50540 55300 50596 55310
rect 50540 55206 50596 55244
rect 51212 55298 51268 55310
rect 51212 55246 51214 55298
rect 51266 55246 51268 55298
rect 49756 55022 49758 55074
rect 49810 55022 49812 55074
rect 49756 54964 49812 55022
rect 50988 55186 51044 55198
rect 50988 55134 50990 55186
rect 51042 55134 51044 55186
rect 50988 54964 51044 55134
rect 49756 54898 49812 54908
rect 50556 54908 50820 54918
rect 49532 54852 49588 54862
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 49532 54626 49588 54796
rect 50988 54740 51044 54908
rect 51212 54964 51268 55246
rect 51212 54898 51268 54908
rect 50764 54684 51044 54740
rect 49532 54574 49534 54626
rect 49586 54574 49588 54626
rect 49532 54562 49588 54574
rect 49644 54628 49700 54638
rect 49644 53956 49700 54572
rect 49868 54516 49924 54526
rect 49868 54422 49924 54460
rect 50204 54516 50260 54526
rect 50204 54422 50260 54460
rect 49644 53862 49700 53900
rect 49980 54402 50036 54414
rect 49980 54350 49982 54402
rect 50034 54350 50036 54402
rect 49420 53678 49422 53730
rect 49474 53678 49476 53730
rect 49420 50596 49476 53678
rect 49756 53844 49812 53854
rect 49756 53730 49812 53788
rect 49756 53678 49758 53730
rect 49810 53678 49812 53730
rect 49644 53508 49700 53518
rect 49532 53506 49700 53508
rect 49532 53454 49646 53506
rect 49698 53454 49700 53506
rect 49532 53452 49700 53454
rect 49532 52386 49588 53452
rect 49644 53442 49700 53452
rect 49756 52946 49812 53678
rect 49756 52894 49758 52946
rect 49810 52894 49812 52946
rect 49756 52882 49812 52894
rect 49532 52334 49534 52386
rect 49586 52334 49588 52386
rect 49532 52322 49588 52334
rect 49868 52722 49924 52734
rect 49868 52670 49870 52722
rect 49922 52670 49924 52722
rect 49644 52164 49700 52174
rect 49644 51604 49700 52108
rect 49644 51510 49700 51548
rect 49420 49140 49476 50540
rect 49756 51268 49812 51278
rect 49756 50370 49812 51212
rect 49756 50318 49758 50370
rect 49810 50318 49812 50370
rect 49756 50036 49812 50318
rect 49644 49980 49812 50036
rect 49532 49698 49588 49710
rect 49532 49646 49534 49698
rect 49586 49646 49588 49698
rect 49532 49588 49588 49646
rect 49532 49522 49588 49532
rect 49308 49028 49364 49038
rect 49420 49028 49476 49084
rect 49532 49028 49588 49038
rect 49420 49026 49588 49028
rect 49420 48974 49534 49026
rect 49586 48974 49588 49026
rect 49420 48972 49588 48974
rect 49308 48934 49364 48972
rect 49532 48962 49588 48972
rect 49644 49028 49700 49980
rect 49644 48934 49700 48972
rect 49756 49812 49812 49822
rect 49196 48412 49700 48468
rect 49644 48354 49700 48412
rect 49644 48302 49646 48354
rect 49698 48302 49700 48354
rect 48748 47740 49140 47796
rect 48412 47460 48468 47470
rect 48412 47458 48580 47460
rect 48412 47406 48414 47458
rect 48466 47406 48580 47458
rect 48412 47404 48580 47406
rect 48412 47394 48468 47404
rect 48412 46562 48468 46574
rect 48412 46510 48414 46562
rect 48466 46510 48468 46562
rect 48412 45668 48468 46510
rect 48412 45602 48468 45612
rect 48524 45890 48580 47404
rect 48748 46898 48804 47740
rect 48748 46846 48750 46898
rect 48802 46846 48804 46898
rect 48748 46834 48804 46846
rect 48972 47570 49028 47582
rect 48972 47518 48974 47570
rect 49026 47518 49028 47570
rect 48972 47012 49028 47518
rect 48524 45838 48526 45890
rect 48578 45838 48580 45890
rect 48524 45332 48580 45838
rect 48972 45668 49028 46956
rect 48972 45602 49028 45612
rect 48636 45332 48692 45342
rect 48524 45276 48636 45332
rect 48636 45200 48692 45276
rect 48300 44492 48580 44548
rect 47852 44034 47908 44044
rect 48076 44100 48132 44110
rect 48076 44006 48132 44044
rect 48300 43428 48356 43438
rect 48300 43334 48356 43372
rect 48188 42756 48244 42766
rect 48188 42662 48244 42700
rect 47740 42532 47796 42542
rect 47740 42438 47796 42476
rect 48300 41860 48356 41870
rect 48300 41766 48356 41804
rect 47516 41188 47572 41198
rect 47516 41186 48132 41188
rect 47516 41134 47518 41186
rect 47570 41134 48132 41186
rect 47516 41132 48132 41134
rect 47516 41122 47572 41132
rect 47628 40964 47684 40974
rect 47404 40292 47460 40302
rect 47404 39730 47460 40236
rect 47404 39678 47406 39730
rect 47458 39678 47460 39730
rect 47404 39508 47460 39678
rect 47404 39442 47460 39452
rect 47180 38612 47348 38668
rect 47180 34244 47236 34254
rect 47180 34150 47236 34188
rect 44940 31892 45332 31948
rect 47068 31892 47236 31948
rect 44828 27748 44884 27758
rect 44716 27746 44884 27748
rect 44716 27694 44830 27746
rect 44882 27694 44884 27746
rect 44716 27692 44884 27694
rect 44716 26964 44772 27692
rect 44828 27682 44884 27692
rect 44716 26870 44772 26908
rect 44716 24610 44772 24622
rect 44716 24558 44718 24610
rect 44770 24558 44772 24610
rect 44716 23828 44772 24558
rect 44716 23734 44772 23772
rect 44268 22148 44324 22158
rect 44268 21586 44324 22092
rect 45052 22036 45108 22046
rect 44492 21700 44548 21710
rect 44492 21606 44548 21644
rect 44268 21534 44270 21586
rect 44322 21534 44324 21586
rect 44268 21522 44324 21534
rect 45052 21476 45108 21980
rect 45052 21382 45108 21420
rect 43596 6626 43652 6636
rect 45276 6356 45332 31892
rect 45500 28532 45556 28542
rect 45500 28530 45780 28532
rect 45500 28478 45502 28530
rect 45554 28478 45780 28530
rect 45500 28476 45780 28478
rect 45500 28466 45556 28476
rect 45724 27298 45780 28476
rect 45836 28420 45892 28430
rect 45836 28418 47012 28420
rect 45836 28366 45838 28418
rect 45890 28366 47012 28418
rect 45836 28364 47012 28366
rect 45836 28354 45892 28364
rect 46956 27970 47012 28364
rect 46956 27918 46958 27970
rect 47010 27918 47012 27970
rect 46956 27906 47012 27918
rect 45724 27246 45726 27298
rect 45778 27246 45780 27298
rect 45724 27234 45780 27246
rect 46060 27300 46116 27310
rect 46060 27206 46116 27244
rect 46844 27188 46900 27198
rect 46844 27074 46900 27132
rect 46844 27022 46846 27074
rect 46898 27022 46900 27074
rect 46844 27010 46900 27022
rect 46620 26964 46676 26974
rect 46620 26870 46676 26908
rect 45612 25506 45668 25518
rect 45612 25454 45614 25506
rect 45666 25454 45668 25506
rect 45612 24164 45668 25454
rect 45836 25284 45892 25294
rect 45836 25282 46900 25284
rect 45836 25230 45838 25282
rect 45890 25230 46900 25282
rect 45836 25228 46900 25230
rect 45836 25218 45892 25228
rect 46844 24834 46900 25228
rect 46844 24782 46846 24834
rect 46898 24782 46900 24834
rect 46844 24770 46900 24782
rect 45724 24164 45780 24174
rect 45612 24162 45780 24164
rect 45612 24110 45726 24162
rect 45778 24110 45780 24162
rect 45612 24108 45780 24110
rect 45724 24098 45780 24108
rect 46060 23940 46116 23950
rect 46060 23846 46116 23884
rect 46844 23938 46900 23950
rect 46844 23886 46846 23938
rect 46898 23886 46900 23938
rect 46620 23828 46676 23838
rect 46620 23734 46676 23772
rect 46844 23716 46900 23886
rect 46844 23650 46900 23660
rect 45836 23266 45892 23278
rect 45836 23214 45838 23266
rect 45890 23214 45892 23266
rect 45612 23154 45668 23166
rect 45612 23102 45614 23154
rect 45666 23102 45668 23154
rect 45500 22146 45556 22158
rect 45500 22094 45502 22146
rect 45554 22094 45556 22146
rect 45500 22036 45556 22094
rect 45500 21970 45556 21980
rect 45500 20914 45556 20926
rect 45500 20862 45502 20914
rect 45554 20862 45556 20914
rect 45500 20132 45556 20862
rect 45612 20188 45668 23102
rect 45836 20916 45892 23214
rect 47180 22484 47236 31892
rect 47292 27300 47348 38612
rect 47292 27188 47348 27244
rect 47404 27188 47460 27198
rect 47292 27186 47460 27188
rect 47292 27134 47406 27186
rect 47458 27134 47460 27186
rect 47292 27132 47460 27134
rect 47404 27122 47460 27132
rect 47628 26068 47684 40908
rect 47740 40964 47796 40974
rect 47740 40962 48020 40964
rect 47740 40910 47742 40962
rect 47794 40910 48020 40962
rect 47740 40908 48020 40910
rect 47740 40898 47796 40908
rect 47964 40514 48020 40908
rect 47964 40462 47966 40514
rect 48018 40462 48020 40514
rect 47964 40450 48020 40462
rect 48076 39842 48132 41132
rect 48076 39790 48078 39842
rect 48130 39790 48132 39842
rect 48076 39778 48132 39790
rect 48412 39732 48468 39742
rect 48412 39638 48468 39676
rect 47964 34130 48020 34142
rect 47964 34078 47966 34130
rect 48018 34078 48020 34130
rect 47964 34020 48020 34078
rect 48412 34020 48468 34030
rect 47964 34018 48468 34020
rect 47964 33966 48414 34018
rect 48466 33966 48468 34018
rect 47964 33964 48468 33966
rect 47740 33460 47796 33470
rect 47740 33366 47796 33404
rect 48188 33348 48244 33358
rect 48188 33254 48244 33292
rect 48188 32004 48244 32014
rect 47740 29426 47796 29438
rect 47740 29374 47742 29426
rect 47794 29374 47796 29426
rect 47740 28532 47796 29374
rect 47740 28466 47796 28476
rect 48188 28082 48244 31948
rect 48412 32004 48468 33964
rect 48524 33460 48580 44492
rect 49084 44546 49140 47740
rect 49532 48242 49588 48254
rect 49532 48190 49534 48242
rect 49586 48190 49588 48242
rect 49532 47012 49588 48190
rect 49532 46946 49588 46956
rect 49196 45668 49252 45678
rect 49196 45574 49252 45612
rect 49644 45666 49700 48302
rect 49644 45614 49646 45666
rect 49698 45614 49700 45666
rect 49420 45332 49476 45342
rect 49420 45238 49476 45276
rect 49084 44494 49086 44546
rect 49138 44494 49140 44546
rect 49084 44434 49140 44494
rect 49084 44382 49086 44434
rect 49138 44382 49140 44434
rect 48860 43426 48916 43438
rect 48860 43374 48862 43426
rect 48914 43374 48916 43426
rect 48860 43092 48916 43374
rect 48860 43026 48916 43036
rect 48748 42868 48804 42878
rect 49084 42868 49140 44382
rect 49532 44098 49588 44110
rect 49532 44046 49534 44098
rect 49586 44046 49588 44098
rect 49532 43652 49588 44046
rect 49532 43586 49588 43596
rect 48748 42866 49140 42868
rect 48748 42814 48750 42866
rect 48802 42814 49140 42866
rect 48748 42812 49140 42814
rect 49532 43428 49588 43438
rect 48748 42802 48804 42812
rect 49532 42754 49588 43372
rect 49532 42702 49534 42754
rect 49586 42702 49588 42754
rect 49532 42690 49588 42702
rect 48972 42642 49028 42654
rect 48972 42590 48974 42642
rect 49026 42590 49028 42642
rect 48748 41858 48804 41870
rect 48748 41806 48750 41858
rect 48802 41806 48804 41858
rect 48748 41748 48804 41806
rect 48748 41682 48804 41692
rect 48972 41300 49028 42590
rect 49196 41300 49252 41310
rect 48972 41298 49252 41300
rect 48972 41246 49198 41298
rect 49250 41246 49252 41298
rect 48972 41244 49252 41246
rect 49196 40964 49252 41244
rect 49196 40898 49252 40908
rect 49420 41188 49476 41198
rect 49420 40626 49476 41132
rect 49420 40574 49422 40626
rect 49474 40574 49476 40626
rect 48748 40404 48804 40414
rect 48748 40310 48804 40348
rect 49420 40404 49476 40574
rect 49420 40338 49476 40348
rect 49644 39732 49700 45614
rect 49756 43204 49812 49756
rect 49868 49588 49924 52670
rect 49980 52388 50036 54350
rect 50204 53730 50260 53742
rect 50204 53678 50206 53730
rect 50258 53678 50260 53730
rect 50092 52388 50148 52398
rect 49980 52386 50148 52388
rect 49980 52334 50094 52386
rect 50146 52334 50148 52386
rect 49980 52332 50148 52334
rect 50092 52322 50148 52332
rect 50204 52276 50260 53678
rect 50652 53732 50708 53742
rect 50540 53620 50596 53630
rect 50540 53526 50596 53564
rect 50652 53508 50708 53676
rect 50764 53620 50820 54684
rect 51212 54516 51268 54526
rect 51212 54422 51268 54460
rect 50876 54404 50932 54414
rect 50876 54310 50932 54348
rect 51324 53956 51380 57708
rect 51436 57538 51492 57550
rect 51436 57486 51438 57538
rect 51490 57486 51492 57538
rect 51436 57204 51492 57486
rect 51436 57138 51492 57148
rect 51436 56644 51492 56654
rect 51548 56644 51604 56654
rect 51436 56642 51548 56644
rect 51436 56590 51438 56642
rect 51490 56590 51548 56642
rect 51436 56588 51548 56590
rect 51436 56578 51492 56588
rect 51436 55970 51492 55982
rect 51436 55918 51438 55970
rect 51490 55918 51492 55970
rect 51436 55748 51492 55918
rect 51548 55860 51604 56588
rect 51548 55794 51604 55804
rect 51436 55300 51492 55692
rect 51548 55300 51604 55310
rect 51436 55298 51604 55300
rect 51436 55246 51550 55298
rect 51602 55246 51604 55298
rect 51436 55244 51604 55246
rect 51436 55074 51492 55086
rect 51436 55022 51438 55074
rect 51490 55022 51492 55074
rect 51436 54626 51492 55022
rect 51436 54574 51438 54626
rect 51490 54574 51492 54626
rect 51436 54562 51492 54574
rect 51548 54740 51604 55244
rect 50764 53554 50820 53564
rect 50876 53900 51380 53956
rect 51436 54292 51492 54302
rect 50652 53442 50708 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50428 52946 50484 52958
rect 50428 52894 50430 52946
rect 50482 52894 50484 52946
rect 50428 52612 50484 52894
rect 50428 52546 50484 52556
rect 50428 52386 50484 52398
rect 50428 52334 50430 52386
rect 50482 52334 50484 52386
rect 50428 52276 50484 52334
rect 50204 52220 50484 52276
rect 49980 51940 50036 51950
rect 49980 51266 50036 51884
rect 49980 51214 49982 51266
rect 50034 51214 50036 51266
rect 49980 49812 50036 51214
rect 50316 51940 50372 51950
rect 50204 50484 50260 50522
rect 50204 50418 50260 50428
rect 49980 49746 50036 49756
rect 50204 49810 50260 49822
rect 50204 49758 50206 49810
rect 50258 49758 50260 49810
rect 49868 49532 50036 49588
rect 49980 49026 50036 49532
rect 49980 48974 49982 49026
rect 50034 48974 50036 49026
rect 49980 48962 50036 48974
rect 50092 49028 50148 49038
rect 49868 48356 49924 48366
rect 49868 48262 49924 48300
rect 49868 46900 49924 46910
rect 49868 46676 49924 46844
rect 49868 46582 49924 46620
rect 49980 46562 50036 46574
rect 49980 46510 49982 46562
rect 50034 46510 50036 46562
rect 49980 45668 50036 46510
rect 50092 46004 50148 48972
rect 50204 48692 50260 49758
rect 50316 49812 50372 51884
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50428 51604 50484 51614
rect 50428 51268 50484 51548
rect 50876 51492 50932 53900
rect 50988 53732 51044 53742
rect 50988 53638 51044 53676
rect 51324 53508 51380 53518
rect 51324 53170 51380 53452
rect 51324 53118 51326 53170
rect 51378 53118 51380 53170
rect 51324 53106 51380 53118
rect 51100 52162 51156 52174
rect 51100 52110 51102 52162
rect 51154 52110 51156 52162
rect 50988 51940 51044 51950
rect 50988 51846 51044 51884
rect 51100 51716 51156 52110
rect 51100 51650 51156 51660
rect 51436 51716 51492 54236
rect 51548 54068 51604 54684
rect 51548 54002 51604 54012
rect 51660 54964 51716 54974
rect 51436 51650 51492 51660
rect 51548 53844 51604 53854
rect 51548 51602 51604 53788
rect 51548 51550 51550 51602
rect 51602 51550 51604 51602
rect 51548 51538 51604 51550
rect 51660 53618 51716 54908
rect 51772 54852 51828 59836
rect 52220 58660 52276 60622
rect 53004 60674 53060 60686
rect 53004 60622 53006 60674
rect 53058 60622 53060 60674
rect 52892 60564 52948 60574
rect 52780 59892 52836 59902
rect 52780 59798 52836 59836
rect 52332 59778 52388 59790
rect 52332 59726 52334 59778
rect 52386 59726 52388 59778
rect 52332 59444 52388 59726
rect 52332 59378 52388 59388
rect 52892 59330 52948 60508
rect 53004 60452 53060 60622
rect 53004 60386 53060 60396
rect 52892 59278 52894 59330
rect 52946 59278 52948 59330
rect 52892 59266 52948 59278
rect 52220 58546 52276 58604
rect 52220 58494 52222 58546
rect 52274 58494 52276 58546
rect 52220 58482 52276 58494
rect 52780 58996 52836 59006
rect 52780 58546 52836 58940
rect 52780 58494 52782 58546
rect 52834 58494 52836 58546
rect 52780 58482 52836 58494
rect 51996 58324 52052 58334
rect 51996 57874 52052 58268
rect 51996 57822 51998 57874
rect 52050 57822 52052 57874
rect 51996 57652 52052 57822
rect 52444 57876 52500 57886
rect 52444 57782 52500 57820
rect 51996 57586 52052 57596
rect 52892 57650 52948 57662
rect 52892 57598 52894 57650
rect 52946 57598 52948 57650
rect 52668 57540 52724 57550
rect 52444 57316 52500 57326
rect 52220 56644 52276 56654
rect 52220 56550 52276 56588
rect 52332 56308 52388 56318
rect 52332 56084 52388 56252
rect 52332 55990 52388 56028
rect 51884 55970 51940 55982
rect 51884 55918 51886 55970
rect 51938 55918 51940 55970
rect 51884 55858 51940 55918
rect 51884 55806 51886 55858
rect 51938 55806 51940 55858
rect 51884 55794 51940 55806
rect 51996 55972 52052 55982
rect 51772 54786 51828 54796
rect 51884 55524 51940 55534
rect 51884 54738 51940 55468
rect 51996 55412 52052 55916
rect 51996 55346 52052 55356
rect 52332 55412 52388 55422
rect 52332 55298 52388 55356
rect 52332 55246 52334 55298
rect 52386 55246 52388 55298
rect 52108 55186 52164 55198
rect 52108 55134 52110 55186
rect 52162 55134 52164 55186
rect 52108 55076 52164 55134
rect 52108 55010 52164 55020
rect 51884 54686 51886 54738
rect 51938 54686 51940 54738
rect 51884 54674 51940 54686
rect 52220 54740 52276 54750
rect 51772 54626 51828 54638
rect 51772 54574 51774 54626
rect 51826 54574 51828 54626
rect 51772 54514 51828 54574
rect 51772 54462 51774 54514
rect 51826 54462 51828 54514
rect 51772 54450 51828 54462
rect 52220 54514 52276 54684
rect 52220 54462 52222 54514
rect 52274 54462 52276 54514
rect 52220 54450 52276 54462
rect 51996 54292 52052 54302
rect 51996 54290 52164 54292
rect 51996 54238 51998 54290
rect 52050 54238 52164 54290
rect 51996 54236 52164 54238
rect 51996 54226 52052 54236
rect 52108 54180 52164 54236
rect 51884 54068 51940 54078
rect 51884 53730 51940 54012
rect 51884 53678 51886 53730
rect 51938 53678 51940 53730
rect 51884 53666 51940 53678
rect 51996 53732 52052 53742
rect 51660 53566 51662 53618
rect 51714 53566 51716 53618
rect 51660 53396 51716 53566
rect 51660 51604 51716 53340
rect 51772 53620 51828 53630
rect 51772 52612 51828 53564
rect 51996 53396 52052 53676
rect 52108 53508 52164 54124
rect 52332 53844 52388 55246
rect 52444 55076 52500 57260
rect 52668 56868 52724 57484
rect 52892 57204 52948 57598
rect 52892 57138 52948 57148
rect 52668 56774 52724 56812
rect 53116 56308 53172 115948
rect 55692 115554 55748 119200
rect 56028 116564 56084 116574
rect 56364 116564 56420 119200
rect 57932 117460 57988 119200
rect 57932 117404 58324 117460
rect 56028 116562 56420 116564
rect 56028 116510 56030 116562
rect 56082 116510 56420 116562
rect 56028 116508 56420 116510
rect 56028 116498 56084 116508
rect 56364 116340 56420 116508
rect 58156 116564 58212 116574
rect 58156 116470 58212 116508
rect 56812 116340 56868 116350
rect 56364 116338 56868 116340
rect 56364 116286 56814 116338
rect 56866 116286 56868 116338
rect 56364 116284 56868 116286
rect 56812 116274 56868 116284
rect 55692 115502 55694 115554
rect 55746 115502 55748 115554
rect 55692 115490 55748 115502
rect 56364 116116 56420 116126
rect 54460 113876 54516 113886
rect 54460 68292 54516 113820
rect 56364 90748 56420 116060
rect 56476 115666 56532 115678
rect 56476 115614 56478 115666
rect 56530 115614 56532 115666
rect 56476 114660 56532 115614
rect 57820 115666 57876 115678
rect 57820 115614 57822 115666
rect 57874 115614 57876 115666
rect 56924 114772 56980 114782
rect 56924 114678 56980 114716
rect 57484 114772 57540 114782
rect 57484 114678 57540 114716
rect 57820 114770 57876 115614
rect 58268 115554 58324 117404
rect 59276 115892 59332 119200
rect 59276 115826 59332 115836
rect 59500 116564 59556 116574
rect 59388 115668 59444 115678
rect 58268 115502 58270 115554
rect 58322 115502 58324 115554
rect 58268 115490 58324 115502
rect 59164 115666 59444 115668
rect 59164 115614 59390 115666
rect 59442 115614 59444 115666
rect 59164 115612 59444 115614
rect 57820 114718 57822 114770
rect 57874 114718 57876 114770
rect 57820 114706 57876 114718
rect 59164 114994 59220 115612
rect 59388 115602 59444 115612
rect 59164 114942 59166 114994
rect 59218 114942 59220 114994
rect 56476 114566 56532 114604
rect 56924 102452 56980 102462
rect 56364 90692 56868 90748
rect 55916 69186 55972 69198
rect 55916 69134 55918 69186
rect 55970 69134 55972 69186
rect 55916 68852 55972 69134
rect 55916 68786 55972 68796
rect 56476 68852 56532 68862
rect 54460 68226 54516 68236
rect 55244 68514 55300 68526
rect 55244 68462 55246 68514
rect 55298 68462 55300 68514
rect 52668 56252 53172 56308
rect 53228 68180 53284 68190
rect 53228 56308 53284 68124
rect 53900 68068 53956 68078
rect 53340 66948 53396 66958
rect 53340 66946 53732 66948
rect 53340 66894 53342 66946
rect 53394 66894 53732 66946
rect 53340 66892 53732 66894
rect 53340 66882 53396 66892
rect 53676 66498 53732 66892
rect 53676 66446 53678 66498
rect 53730 66446 53732 66498
rect 53676 66434 53732 66446
rect 53788 66050 53844 66062
rect 53788 65998 53790 66050
rect 53842 65998 53844 66050
rect 53788 65604 53844 65998
rect 53676 65548 53844 65604
rect 53340 65492 53396 65502
rect 53340 65398 53396 65436
rect 53676 64484 53732 65548
rect 53900 65492 53956 68012
rect 54908 67954 54964 67966
rect 54908 67902 54910 67954
rect 54962 67902 54964 67954
rect 54908 67172 54964 67902
rect 54908 67106 54964 67116
rect 55132 67842 55188 67854
rect 55132 67790 55134 67842
rect 55186 67790 55188 67842
rect 54796 66500 54852 66510
rect 54236 66276 54292 66286
rect 54012 66164 54068 66174
rect 54012 66070 54068 66108
rect 53900 65426 53956 65436
rect 53452 64428 53676 64484
rect 53452 64146 53508 64428
rect 53676 64418 53732 64428
rect 53788 65378 53844 65390
rect 53788 65326 53790 65378
rect 53842 65326 53844 65378
rect 53788 64260 53844 65326
rect 54236 65378 54292 66220
rect 54572 66274 54628 66286
rect 54572 66222 54574 66274
rect 54626 66222 54628 66274
rect 54572 65492 54628 66222
rect 54796 66274 54852 66444
rect 54796 66222 54798 66274
rect 54850 66222 54852 66274
rect 54684 65940 54740 65950
rect 54684 65714 54740 65884
rect 54684 65662 54686 65714
rect 54738 65662 54740 65714
rect 54684 65650 54740 65662
rect 54796 65716 54852 66222
rect 54908 66274 54964 66286
rect 54908 66222 54910 66274
rect 54962 66222 54964 66274
rect 54908 65940 54964 66222
rect 54908 65874 54964 65884
rect 55020 65716 55076 65726
rect 54796 65714 55076 65716
rect 54796 65662 55022 65714
rect 55074 65662 55076 65714
rect 54796 65660 55076 65662
rect 54572 65426 54628 65436
rect 54236 65326 54238 65378
rect 54290 65326 54292 65378
rect 54236 65156 54292 65326
rect 54236 65090 54292 65100
rect 54236 64484 54292 64494
rect 54292 64428 54404 64484
rect 54236 64352 54292 64428
rect 54012 64260 54068 64270
rect 53788 64204 54012 64260
rect 53452 64094 53454 64146
rect 53506 64094 53508 64146
rect 53452 64082 53508 64094
rect 53452 63364 53508 63374
rect 53340 62244 53396 62282
rect 53340 62178 53396 62188
rect 53452 62188 53508 63308
rect 53564 63138 53620 63150
rect 53564 63086 53566 63138
rect 53618 63086 53620 63138
rect 53564 62580 53620 63086
rect 53564 62514 53620 62524
rect 53788 62242 53844 62254
rect 53788 62190 53790 62242
rect 53842 62190 53844 62242
rect 53788 62188 53844 62190
rect 53452 62132 53844 62188
rect 53564 61682 53620 62132
rect 53900 62130 53956 62142
rect 53900 62078 53902 62130
rect 53954 62078 53956 62130
rect 53564 61630 53566 61682
rect 53618 61630 53620 61682
rect 53564 61618 53620 61630
rect 53788 61796 53844 61806
rect 53676 61236 53732 61246
rect 53564 60788 53620 60798
rect 53564 60694 53620 60732
rect 53564 60004 53620 60014
rect 53676 60004 53732 61180
rect 53788 61012 53844 61740
rect 53900 61572 53956 62078
rect 54012 61794 54068 64204
rect 54012 61742 54014 61794
rect 54066 61742 54068 61794
rect 54012 61730 54068 61742
rect 54124 64148 54180 64158
rect 54348 64148 54404 64428
rect 54124 64146 54404 64148
rect 54124 64094 54126 64146
rect 54178 64094 54404 64146
rect 54124 64092 54404 64094
rect 54124 61796 54180 64092
rect 54348 63924 54404 64092
rect 54348 63858 54404 63868
rect 54236 63810 54292 63822
rect 54236 63758 54238 63810
rect 54290 63758 54292 63810
rect 54236 63250 54292 63758
rect 54348 63700 54404 63710
rect 54348 63606 54404 63644
rect 54236 63198 54238 63250
rect 54290 63198 54292 63250
rect 54236 63186 54292 63198
rect 54684 62580 54740 62590
rect 54796 62580 54852 65660
rect 55020 65650 55076 65660
rect 55132 65716 55188 67790
rect 55244 67060 55300 68462
rect 55692 68516 55748 68526
rect 55692 68514 55860 68516
rect 55692 68462 55694 68514
rect 55746 68462 55860 68514
rect 55692 68460 55860 68462
rect 55692 68450 55748 68460
rect 55692 67732 55748 67742
rect 55580 67730 55748 67732
rect 55580 67678 55694 67730
rect 55746 67678 55748 67730
rect 55580 67676 55748 67678
rect 55580 67284 55636 67676
rect 55692 67666 55748 67676
rect 55244 66994 55300 67004
rect 55356 67228 55636 67284
rect 55356 66836 55412 67228
rect 55692 67172 55748 67182
rect 55580 66948 55636 66958
rect 55580 66854 55636 66892
rect 55244 66780 55412 66836
rect 55244 66274 55300 66780
rect 55244 66222 55246 66274
rect 55298 66222 55300 66274
rect 55244 66210 55300 66222
rect 55468 66386 55524 66398
rect 55468 66334 55470 66386
rect 55522 66334 55524 66386
rect 55356 66164 55412 66174
rect 55356 66050 55412 66108
rect 55356 65998 55358 66050
rect 55410 65998 55412 66050
rect 55356 65986 55412 65998
rect 54908 64820 54964 64830
rect 55132 64820 55188 65660
rect 55468 64932 55524 66334
rect 55580 65716 55636 65726
rect 55692 65716 55748 67116
rect 55804 66052 55860 68460
rect 56140 68514 56196 68526
rect 56140 68462 56142 68514
rect 56194 68462 56196 68514
rect 56140 66500 56196 68462
rect 56476 68514 56532 68796
rect 56476 68462 56478 68514
rect 56530 68462 56532 68514
rect 56252 67172 56308 67182
rect 56252 67078 56308 67116
rect 56364 67172 56420 67182
rect 56476 67172 56532 68462
rect 56588 67954 56644 67966
rect 56588 67902 56590 67954
rect 56642 67902 56644 67954
rect 56588 67282 56644 67902
rect 56700 67842 56756 67854
rect 56700 67790 56702 67842
rect 56754 67790 56756 67842
rect 56700 67620 56756 67790
rect 56700 67554 56756 67564
rect 56588 67230 56590 67282
rect 56642 67230 56644 67282
rect 56588 67218 56644 67230
rect 56364 67170 56532 67172
rect 56364 67118 56366 67170
rect 56418 67118 56532 67170
rect 56364 67116 56532 67118
rect 56140 66434 56196 66444
rect 56364 66948 56420 67116
rect 55916 66388 55972 66398
rect 55916 66294 55972 66332
rect 55804 65986 55860 65996
rect 55580 65714 55748 65716
rect 55580 65662 55582 65714
rect 55634 65662 55748 65714
rect 55580 65660 55748 65662
rect 56364 65716 56420 66892
rect 56588 66500 56644 66510
rect 56588 66274 56644 66444
rect 56588 66222 56590 66274
rect 56642 66222 56644 66274
rect 56588 66210 56644 66222
rect 56700 66274 56756 66286
rect 56700 66222 56702 66274
rect 56754 66222 56756 66274
rect 56476 66052 56532 66062
rect 56476 65958 56532 65996
rect 55580 65650 55636 65660
rect 56364 65650 56420 65660
rect 56700 65940 56756 66222
rect 54908 64818 55188 64820
rect 54908 64766 54910 64818
rect 54962 64766 55188 64818
rect 54908 64764 55188 64766
rect 55244 64876 55524 64932
rect 55916 65380 55972 65390
rect 54908 64754 54964 64764
rect 55244 64260 55300 64876
rect 55356 64708 55412 64718
rect 55356 64614 55412 64652
rect 55916 64708 55972 65324
rect 55692 64484 55748 64494
rect 55244 64194 55300 64204
rect 55356 64482 55748 64484
rect 55356 64430 55694 64482
rect 55746 64430 55748 64482
rect 55356 64428 55748 64430
rect 55356 63922 55412 64428
rect 55692 64418 55748 64428
rect 55356 63870 55358 63922
rect 55410 63870 55412 63922
rect 54908 63812 54964 63822
rect 54908 63810 55188 63812
rect 54908 63758 54910 63810
rect 54962 63758 55188 63810
rect 54908 63756 55188 63758
rect 54908 63746 54964 63756
rect 54684 62578 54852 62580
rect 54684 62526 54686 62578
rect 54738 62526 54852 62578
rect 54684 62524 54852 62526
rect 54684 62514 54740 62524
rect 54796 62468 54852 62524
rect 54796 62402 54852 62412
rect 55132 62466 55188 63756
rect 55244 63700 55300 63710
rect 55244 62578 55300 63644
rect 55356 63588 55412 63870
rect 55804 63924 55860 63934
rect 55916 63924 55972 64652
rect 55804 63922 55972 63924
rect 55804 63870 55806 63922
rect 55858 63870 55972 63922
rect 55804 63868 55972 63870
rect 56140 65380 56196 65390
rect 56588 65380 56644 65390
rect 56140 65378 56644 65380
rect 56140 65326 56142 65378
rect 56194 65326 56590 65378
rect 56642 65326 56644 65378
rect 56140 65324 56644 65326
rect 56140 64708 56196 65324
rect 56588 65314 56644 65324
rect 56700 65156 56756 65884
rect 56700 65090 56756 65100
rect 55804 63858 55860 63868
rect 55356 63522 55412 63532
rect 56140 63588 56196 64652
rect 56700 64148 56756 64158
rect 56812 64148 56868 90692
rect 56700 64146 56812 64148
rect 56700 64094 56702 64146
rect 56754 64094 56812 64146
rect 56700 64092 56812 64094
rect 56700 64082 56756 64092
rect 56812 64016 56868 64092
rect 56140 63522 56196 63532
rect 56364 63588 56420 63598
rect 56364 63250 56420 63532
rect 56364 63198 56366 63250
rect 56418 63198 56420 63250
rect 56364 63186 56420 63198
rect 55244 62526 55246 62578
rect 55298 62526 55300 62578
rect 55244 62514 55300 62526
rect 55916 63140 55972 63150
rect 56924 63140 56980 102396
rect 57932 93044 57988 93054
rect 57036 68066 57092 68078
rect 57036 68014 57038 68066
rect 57090 68014 57092 68066
rect 57036 66274 57092 68014
rect 57820 67620 57876 67630
rect 57820 67526 57876 67564
rect 57596 67060 57652 67070
rect 57596 66966 57652 67004
rect 57036 66222 57038 66274
rect 57090 66222 57092 66274
rect 57036 66210 57092 66222
rect 57260 66386 57316 66398
rect 57260 66334 57262 66386
rect 57314 66334 57316 66386
rect 57260 65604 57316 66334
rect 57596 66276 57652 66286
rect 57596 66182 57652 66220
rect 57932 66276 57988 92988
rect 58828 89682 58884 89694
rect 58828 89630 58830 89682
rect 58882 89630 58884 89682
rect 58828 89572 58884 89630
rect 59164 89682 59220 114942
rect 59500 102508 59556 116508
rect 59948 116564 60004 116574
rect 59948 116470 60004 116508
rect 60508 116564 60564 119200
rect 60508 116498 60564 116508
rect 60956 116564 61012 116574
rect 61740 116564 61796 116574
rect 60956 116562 61124 116564
rect 60956 116510 60958 116562
rect 61010 116510 61124 116562
rect 60956 116508 61124 116510
rect 60956 116498 61012 116508
rect 60060 115892 60116 115902
rect 60060 115554 60116 115836
rect 60060 115502 60062 115554
rect 60114 115502 60116 115554
rect 60060 115490 60116 115502
rect 59164 89630 59166 89682
rect 59218 89630 59220 89682
rect 59164 89618 59220 89630
rect 59388 102452 59556 102508
rect 58828 89506 58884 89516
rect 59276 68292 59332 68302
rect 58940 67172 58996 67182
rect 58268 66946 58324 66958
rect 58268 66894 58270 66946
rect 58322 66894 58324 66946
rect 58268 66386 58324 66894
rect 58940 66500 58996 67116
rect 58268 66334 58270 66386
rect 58322 66334 58324 66386
rect 58268 66322 58324 66334
rect 58492 66444 58996 66500
rect 57932 66210 57988 66220
rect 58492 66274 58548 66444
rect 58492 66222 58494 66274
rect 58546 66222 58548 66274
rect 58492 66210 58548 66222
rect 58156 66162 58212 66174
rect 58156 66110 58158 66162
rect 58210 66110 58212 66162
rect 57708 66052 57764 66062
rect 58156 66052 58212 66110
rect 57708 66050 58212 66052
rect 57708 65998 57710 66050
rect 57762 65998 58212 66050
rect 57708 65996 58212 65998
rect 57708 65986 57764 65996
rect 58492 65604 58548 65614
rect 57260 65602 58548 65604
rect 57260 65550 58494 65602
rect 58546 65550 58548 65602
rect 57260 65548 58548 65550
rect 55132 62414 55134 62466
rect 55186 62414 55188 62466
rect 55132 62402 55188 62414
rect 54460 62356 54516 62366
rect 54460 62262 54516 62300
rect 55020 62356 55076 62366
rect 55020 62262 55076 62300
rect 55916 62356 55972 63084
rect 56588 63084 56980 63140
rect 57148 64818 57204 64830
rect 57148 64766 57150 64818
rect 57202 64766 57204 64818
rect 56252 62580 56308 62590
rect 56252 62486 56308 62524
rect 54124 61730 54180 61740
rect 55244 62244 55300 62254
rect 53900 61516 54292 61572
rect 54124 61348 54180 61358
rect 54124 61254 54180 61292
rect 53788 60788 53844 60956
rect 54012 60788 54068 60798
rect 53788 60786 54068 60788
rect 53788 60734 54014 60786
rect 54066 60734 54068 60786
rect 53788 60732 54068 60734
rect 54236 60788 54292 61516
rect 54348 61458 54404 61470
rect 54348 61406 54350 61458
rect 54402 61406 54404 61458
rect 54348 61236 54404 61406
rect 54348 61170 54404 61180
rect 55020 61346 55076 61358
rect 55020 61294 55022 61346
rect 55074 61294 55076 61346
rect 55020 61236 55076 61294
rect 55020 61012 55076 61180
rect 55020 60946 55076 60956
rect 55132 60788 55188 60798
rect 54236 60786 55188 60788
rect 54236 60734 55134 60786
rect 55186 60734 55188 60786
rect 54236 60732 55188 60734
rect 54012 60722 54068 60732
rect 55132 60722 55188 60732
rect 54012 60564 54068 60574
rect 54012 60470 54068 60508
rect 54348 60562 54404 60574
rect 54348 60510 54350 60562
rect 54402 60510 54404 60562
rect 53900 60452 53956 60462
rect 53900 60114 53956 60396
rect 53900 60062 53902 60114
rect 53954 60062 53956 60114
rect 53900 60050 53956 60062
rect 53620 59948 53732 60004
rect 53564 59872 53620 59948
rect 53564 59218 53620 59230
rect 53564 59166 53566 59218
rect 53618 59166 53620 59218
rect 53452 58324 53508 58334
rect 53340 58322 53508 58324
rect 53340 58270 53454 58322
rect 53506 58270 53508 58322
rect 53340 58268 53508 58270
rect 53340 56644 53396 58268
rect 53452 58258 53508 58268
rect 53452 57538 53508 57550
rect 53452 57486 53454 57538
rect 53506 57486 53508 57538
rect 53452 56644 53508 57486
rect 53564 56868 53620 59166
rect 53564 56802 53620 56812
rect 53676 56644 53732 59948
rect 54348 59780 54404 60510
rect 55020 60562 55076 60574
rect 55020 60510 55022 60562
rect 55074 60510 55076 60562
rect 55020 60452 55076 60510
rect 55020 60386 55076 60396
rect 55020 60004 55076 60014
rect 54908 59890 54964 59902
rect 54908 59838 54910 59890
rect 54962 59838 54964 59890
rect 54796 59780 54852 59790
rect 54348 59778 54852 59780
rect 54348 59726 54798 59778
rect 54850 59726 54852 59778
rect 54348 59724 54852 59726
rect 54796 59714 54852 59724
rect 54908 59444 54964 59838
rect 54908 59378 54964 59388
rect 55020 59442 55076 59948
rect 55132 60002 55188 60014
rect 55132 59950 55134 60002
rect 55186 59950 55188 60002
rect 55132 59892 55188 59950
rect 55132 59826 55188 59836
rect 55244 59444 55300 62188
rect 55468 62244 55524 62282
rect 55468 62178 55524 62188
rect 55804 62242 55860 62254
rect 55804 62190 55806 62242
rect 55858 62190 55860 62242
rect 55580 62132 55636 62142
rect 55580 61682 55636 62076
rect 55580 61630 55582 61682
rect 55634 61630 55636 61682
rect 55356 60788 55412 60798
rect 55580 60788 55636 61630
rect 55804 61236 55860 62190
rect 55916 61794 55972 62300
rect 55916 61742 55918 61794
rect 55970 61742 55972 61794
rect 55916 61682 55972 61742
rect 55916 61630 55918 61682
rect 55970 61630 55972 61682
rect 55916 61618 55972 61630
rect 56140 62020 56196 62030
rect 55804 61170 55860 61180
rect 56028 60788 56084 60798
rect 55580 60786 56084 60788
rect 55580 60734 56030 60786
rect 56082 60734 56084 60786
rect 55580 60732 56084 60734
rect 55356 60564 55412 60732
rect 56028 60722 56084 60732
rect 56140 60788 56196 61964
rect 56476 61794 56532 61806
rect 56476 61742 56478 61794
rect 56530 61742 56532 61794
rect 56364 61346 56420 61358
rect 56364 61294 56366 61346
rect 56418 61294 56420 61346
rect 56364 61236 56420 61294
rect 56364 61170 56420 61180
rect 56364 61012 56420 61022
rect 56364 60898 56420 60956
rect 56364 60846 56366 60898
rect 56418 60846 56420 60898
rect 56364 60834 56420 60846
rect 55356 60470 55412 60508
rect 55468 60562 55524 60574
rect 56028 60564 56084 60574
rect 55468 60510 55470 60562
rect 55522 60510 55524 60562
rect 55468 60340 55524 60510
rect 55356 60284 55524 60340
rect 55692 60562 56084 60564
rect 55692 60510 56030 60562
rect 56082 60510 56084 60562
rect 55692 60508 56084 60510
rect 55356 60226 55412 60284
rect 55356 60174 55358 60226
rect 55410 60174 55412 60226
rect 55356 60162 55412 60174
rect 55580 60004 55636 60014
rect 55580 59910 55636 59948
rect 55020 59390 55022 59442
rect 55074 59390 55076 59442
rect 55020 59378 55076 59390
rect 55132 59388 55300 59444
rect 55468 59892 55524 59902
rect 54460 59106 54516 59118
rect 54460 59054 54462 59106
rect 54514 59054 54516 59106
rect 54460 58660 54516 59054
rect 54684 58996 54740 59006
rect 54684 58902 54740 58940
rect 54460 58594 54516 58604
rect 54572 58772 54628 58782
rect 54572 58658 54628 58716
rect 54572 58606 54574 58658
rect 54626 58606 54628 58658
rect 54572 58594 54628 58606
rect 53788 58548 53844 58558
rect 53788 58322 53844 58492
rect 53788 58270 53790 58322
rect 53842 58270 53844 58322
rect 53788 58258 53844 58270
rect 54460 58324 54516 58334
rect 54460 58230 54516 58268
rect 54572 58210 54628 58222
rect 54572 58158 54574 58210
rect 54626 58158 54628 58210
rect 54236 57876 54292 57886
rect 53900 56868 53956 56878
rect 53956 56812 54068 56868
rect 53900 56736 53956 56812
rect 53452 56588 53732 56644
rect 53340 56578 53396 56588
rect 53228 56252 53396 56308
rect 52556 55412 52612 55422
rect 52556 55318 52612 55356
rect 52444 55010 52500 55020
rect 52332 53778 52388 53788
rect 52332 53508 52388 53518
rect 52108 53506 52500 53508
rect 52108 53454 52334 53506
rect 52386 53454 52500 53506
rect 52108 53452 52500 53454
rect 52332 53442 52388 53452
rect 51996 53340 52164 53396
rect 51884 53060 51940 53070
rect 51884 52966 51940 53004
rect 51772 52546 51828 52556
rect 51660 51538 51716 51548
rect 51996 52500 52052 52510
rect 51996 52274 52052 52444
rect 51996 52222 51998 52274
rect 52050 52222 52052 52274
rect 50876 51378 50932 51436
rect 50876 51326 50878 51378
rect 50930 51326 50932 51378
rect 50876 51314 50932 51326
rect 51436 51492 51492 51502
rect 51436 51380 51492 51436
rect 51436 51324 51604 51380
rect 50428 51202 50484 51212
rect 50540 51156 50596 51166
rect 50540 51062 50596 51100
rect 50876 51154 50932 51166
rect 51436 51156 51492 51166
rect 50876 51102 50878 51154
rect 50930 51102 50932 51154
rect 50876 51044 50932 51102
rect 50876 50978 50932 50988
rect 50988 51154 51492 51156
rect 50988 51102 51438 51154
rect 51490 51102 51492 51154
rect 50988 51100 51492 51102
rect 50988 50820 51044 51100
rect 51436 51090 51492 51100
rect 50428 50764 51044 50820
rect 50428 50706 50484 50764
rect 51548 50708 51604 51324
rect 50428 50654 50430 50706
rect 50482 50654 50484 50706
rect 50428 50642 50484 50654
rect 51436 50652 51604 50708
rect 51772 51154 51828 51166
rect 51772 51102 51774 51154
rect 51826 51102 51828 51154
rect 50652 50594 50708 50606
rect 50652 50542 50654 50594
rect 50706 50542 50708 50594
rect 50652 50428 50708 50542
rect 50876 50596 50932 50606
rect 50876 50502 50932 50540
rect 51212 50596 51268 50606
rect 51212 50502 51268 50540
rect 50428 50372 50708 50428
rect 50764 50372 50820 50382
rect 50428 50034 50484 50372
rect 50764 50370 51156 50372
rect 50764 50318 50766 50370
rect 50818 50318 51156 50370
rect 50764 50316 51156 50318
rect 50764 50306 50820 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50988 50148 51044 50158
rect 50428 49982 50430 50034
rect 50482 49982 50484 50034
rect 50428 49970 50484 49982
rect 50876 49924 50932 49934
rect 50988 49924 51044 50092
rect 50876 49922 51044 49924
rect 50876 49870 50878 49922
rect 50930 49870 51044 49922
rect 50876 49868 51044 49870
rect 50876 49858 50932 49868
rect 50428 49812 50484 49822
rect 50316 49810 50484 49812
rect 50316 49758 50430 49810
rect 50482 49758 50484 49810
rect 50316 49756 50484 49758
rect 50428 49746 50484 49756
rect 50540 49810 50596 49822
rect 50540 49758 50542 49810
rect 50594 49758 50596 49810
rect 50540 49252 50596 49758
rect 50428 49196 50596 49252
rect 51100 49250 51156 50316
rect 51100 49198 51102 49250
rect 51154 49198 51156 49250
rect 50316 49140 50372 49150
rect 50316 49046 50372 49084
rect 50204 48132 50260 48636
rect 50204 48066 50260 48076
rect 50316 48802 50372 48814
rect 50316 48750 50318 48802
rect 50370 48750 50372 48802
rect 50316 46116 50372 48750
rect 50428 46900 50484 49196
rect 51100 49186 51156 49198
rect 51324 49364 51380 49374
rect 50540 49026 50596 49038
rect 50540 48974 50542 49026
rect 50594 48974 50596 49026
rect 50540 48916 50596 48974
rect 50540 48850 50596 48860
rect 51212 48802 51268 48814
rect 51212 48750 51214 48802
rect 51266 48750 51268 48802
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50764 48132 50820 48142
rect 50764 48038 50820 48076
rect 51100 47572 51156 47582
rect 51212 47572 51268 48750
rect 51100 47570 51268 47572
rect 51100 47518 51102 47570
rect 51154 47518 51268 47570
rect 51100 47516 51268 47518
rect 51324 48802 51380 49308
rect 51324 48750 51326 48802
rect 51378 48750 51380 48802
rect 51100 47506 51156 47516
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50428 46834 50484 46844
rect 51324 46788 51380 48750
rect 51436 48356 51492 50652
rect 51660 50482 51716 50494
rect 51660 50430 51662 50482
rect 51714 50430 51716 50482
rect 51548 50370 51604 50382
rect 51548 50318 51550 50370
rect 51602 50318 51604 50370
rect 51548 50148 51604 50318
rect 51548 50082 51604 50092
rect 51660 50372 51716 50430
rect 51548 49700 51604 49710
rect 51548 49606 51604 49644
rect 51660 49252 51716 50316
rect 51772 50260 51828 51102
rect 51772 50194 51828 50204
rect 51884 50482 51940 50494
rect 51884 50430 51886 50482
rect 51938 50430 51940 50482
rect 51884 49812 51940 50430
rect 51884 49746 51940 49756
rect 51660 49186 51716 49196
rect 51996 49028 52052 52222
rect 52108 49924 52164 53340
rect 52332 52834 52388 52846
rect 52332 52782 52334 52834
rect 52386 52782 52388 52834
rect 52220 52724 52276 52734
rect 52220 52388 52276 52668
rect 52332 52722 52388 52782
rect 52332 52670 52334 52722
rect 52386 52670 52388 52722
rect 52332 52658 52388 52670
rect 52220 52256 52276 52332
rect 52444 51716 52500 53452
rect 52668 53284 52724 56252
rect 52780 56140 53060 56196
rect 52780 55298 52836 56140
rect 53004 56084 53060 56140
rect 53340 56084 53396 56252
rect 53004 56028 53396 56084
rect 52892 55970 52948 55982
rect 52892 55918 52894 55970
rect 52946 55918 52948 55970
rect 52892 55860 52948 55918
rect 52892 55794 52948 55804
rect 53116 55858 53172 55870
rect 53452 55860 53508 55870
rect 53116 55806 53118 55858
rect 53170 55806 53172 55858
rect 53116 55524 53172 55806
rect 53116 55458 53172 55468
rect 53228 55858 53508 55860
rect 53228 55806 53454 55858
rect 53506 55806 53508 55858
rect 53228 55804 53508 55806
rect 52780 55246 52782 55298
rect 52834 55246 52836 55298
rect 52780 53732 52836 55246
rect 53228 54852 53284 55804
rect 53452 55794 53508 55804
rect 53004 54796 53284 54852
rect 53452 55636 53508 55646
rect 53452 55186 53508 55580
rect 53452 55134 53454 55186
rect 53506 55134 53508 55186
rect 53004 54740 53060 54796
rect 53004 54608 53060 54684
rect 52780 53666 52836 53676
rect 52892 54402 52948 54414
rect 52892 54350 52894 54402
rect 52946 54350 52948 54402
rect 52892 53508 52948 54350
rect 53116 54068 53172 54078
rect 53452 54068 53508 55134
rect 52948 53452 53060 53508
rect 52892 53442 52948 53452
rect 52668 53218 52724 53228
rect 52780 52834 52836 52846
rect 52780 52782 52782 52834
rect 52834 52782 52836 52834
rect 52780 52724 52836 52782
rect 52780 52658 52836 52668
rect 53004 52500 53060 53452
rect 52556 51940 52612 51950
rect 52556 51938 52948 51940
rect 52556 51886 52558 51938
rect 52610 51886 52948 51938
rect 52556 51884 52948 51886
rect 52556 51874 52612 51884
rect 52444 51660 52612 51716
rect 52444 51156 52500 51166
rect 52444 51062 52500 51100
rect 52220 51044 52276 51054
rect 52220 50594 52276 50988
rect 52220 50542 52222 50594
rect 52274 50542 52276 50594
rect 52220 50530 52276 50542
rect 52108 49858 52164 49868
rect 52332 50260 52388 50270
rect 52332 49922 52388 50204
rect 52332 49870 52334 49922
rect 52386 49870 52388 49922
rect 52332 49858 52388 49870
rect 52108 49698 52164 49710
rect 52108 49646 52110 49698
rect 52162 49646 52164 49698
rect 52108 49140 52164 49646
rect 52108 49074 52164 49084
rect 52220 49252 52276 49262
rect 51884 48972 52052 49028
rect 51548 48356 51604 48366
rect 51436 48354 51604 48356
rect 51436 48302 51550 48354
rect 51602 48302 51604 48354
rect 51436 48300 51604 48302
rect 51548 48290 51604 48300
rect 51772 47458 51828 47470
rect 51772 47406 51774 47458
rect 51826 47406 51828 47458
rect 51324 46732 51492 46788
rect 50540 46676 50596 46686
rect 50316 46050 50372 46060
rect 50428 46674 50596 46676
rect 50428 46622 50542 46674
rect 50594 46622 50596 46674
rect 50428 46620 50596 46622
rect 50204 46004 50260 46014
rect 50092 46002 50260 46004
rect 50092 45950 50206 46002
rect 50258 45950 50260 46002
rect 50092 45948 50260 45950
rect 50204 45938 50260 45948
rect 49980 45602 50036 45612
rect 50204 45668 50260 45678
rect 49980 44324 50036 44334
rect 49980 44230 50036 44268
rect 50204 43540 50260 45612
rect 50428 45332 50484 46620
rect 50540 46610 50596 46620
rect 51324 46564 51380 46574
rect 50876 46562 51380 46564
rect 50876 46510 51326 46562
rect 51378 46510 51380 46562
rect 50876 46508 51380 46510
rect 50652 46116 50708 46126
rect 50652 46022 50708 46060
rect 50876 46002 50932 46508
rect 51324 46498 51380 46508
rect 50876 45950 50878 46002
rect 50930 45950 50932 46002
rect 50876 45938 50932 45950
rect 50876 45780 50932 45790
rect 50876 45666 50932 45724
rect 51436 45780 51492 46732
rect 51436 45714 51492 45724
rect 50876 45614 50878 45666
rect 50930 45614 50932 45666
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50428 45266 50484 45276
rect 50540 44994 50596 45006
rect 50540 44942 50542 44994
rect 50594 44942 50596 44994
rect 50540 44660 50596 44942
rect 50540 44594 50596 44604
rect 50876 44660 50932 45614
rect 51548 45666 51604 45678
rect 51548 45614 51550 45666
rect 51602 45614 51604 45666
rect 51548 45556 51604 45614
rect 51548 45490 51604 45500
rect 50988 45332 51044 45342
rect 50988 45238 51044 45276
rect 51436 45332 51492 45342
rect 51436 45238 51492 45276
rect 51772 45332 51828 47406
rect 51772 45266 51828 45276
rect 50932 44604 51044 44660
rect 50876 44594 50932 44604
rect 50316 44546 50372 44558
rect 50316 44494 50318 44546
rect 50370 44494 50372 44546
rect 50316 43652 50372 44494
rect 50428 44436 50484 44446
rect 50428 44342 50484 44380
rect 50876 44100 50932 44110
rect 50876 44006 50932 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50764 43652 50820 43662
rect 50316 43596 50484 43652
rect 50204 43484 50372 43540
rect 49868 43428 49924 43438
rect 49868 43426 50260 43428
rect 49868 43374 49870 43426
rect 49922 43374 50260 43426
rect 49868 43372 50260 43374
rect 49868 43362 49924 43372
rect 49756 43148 50036 43204
rect 49868 42756 49924 42766
rect 49868 42662 49924 42700
rect 49756 42644 49812 42654
rect 49756 42550 49812 42588
rect 49868 41860 49924 41870
rect 49868 41188 49924 41804
rect 49868 41056 49924 41132
rect 49644 39666 49700 39676
rect 49868 39732 49924 39742
rect 49868 39638 49924 39676
rect 49196 39618 49252 39630
rect 49196 39566 49198 39618
rect 49250 39566 49252 39618
rect 48972 39508 49028 39518
rect 48972 39414 49028 39452
rect 49196 39508 49252 39566
rect 48524 33394 48580 33404
rect 48412 31938 48468 31948
rect 48524 33236 48580 33246
rect 48524 29202 48580 33180
rect 49196 31948 49252 39452
rect 49980 31948 50036 43148
rect 50204 42754 50260 43372
rect 50204 42702 50206 42754
rect 50258 42702 50260 42754
rect 50204 42690 50260 42702
rect 50204 39508 50260 39518
rect 50204 39414 50260 39452
rect 49196 31892 49476 31948
rect 48524 29150 48526 29202
rect 48578 29150 48580 29202
rect 48188 28030 48190 28082
rect 48242 28030 48244 28082
rect 47740 27858 47796 27870
rect 47740 27806 47742 27858
rect 47794 27806 47796 27858
rect 47740 27748 47796 27806
rect 48188 27748 48244 28030
rect 47740 27692 48244 27748
rect 48300 28532 48356 28542
rect 47852 27188 47908 27198
rect 47852 27094 47908 27132
rect 47516 26012 47684 26068
rect 47404 23828 47460 23838
rect 47404 23734 47460 23772
rect 46396 22370 46452 22382
rect 46396 22318 46398 22370
rect 46450 22318 46452 22370
rect 46396 22260 46452 22318
rect 47180 22370 47236 22428
rect 47180 22318 47182 22370
rect 47234 22318 47236 22370
rect 47180 22306 47236 22318
rect 46396 22194 46452 22204
rect 46844 22260 46900 22270
rect 46060 22148 46116 22158
rect 46060 22054 46116 22092
rect 45836 20850 45892 20860
rect 45612 20132 46116 20188
rect 45500 20038 45556 20076
rect 46060 20130 46116 20132
rect 46060 20078 46062 20130
rect 46114 20078 46116 20130
rect 46060 20066 46116 20078
rect 46620 20132 46676 20142
rect 46396 19796 46452 19806
rect 46396 19702 46452 19740
rect 46060 6692 46116 6702
rect 45276 6300 45444 6356
rect 43260 5236 43316 5246
rect 43260 5142 43316 5180
rect 43708 4898 43764 4910
rect 43708 4846 43710 4898
rect 43762 4846 43764 4898
rect 43148 4620 43316 4676
rect 43148 4340 43204 4350
rect 42700 4338 43204 4340
rect 42700 4286 43150 4338
rect 43202 4286 43204 4338
rect 42700 4284 43204 4286
rect 43148 4274 43204 4284
rect 42252 4226 42308 4238
rect 42252 4174 42254 4226
rect 42306 4174 42308 4226
rect 41468 3444 41524 3454
rect 42028 3444 42084 3454
rect 41468 3442 42084 3444
rect 41468 3390 41470 3442
rect 41522 3390 42030 3442
rect 42082 3390 42084 3442
rect 41468 3388 42084 3390
rect 41468 3378 41524 3388
rect 30856 200 31080 728
rect 32200 200 32424 728
rect 32508 700 33236 756
rect 33544 200 33768 800
rect 34216 200 34440 800
rect 35532 728 35784 800
rect 35560 200 35784 728
rect 36904 728 37156 800
rect 37576 728 37828 800
rect 36904 200 37128 728
rect 37576 200 37800 728
rect 38920 200 39144 800
rect 40264 728 40516 800
rect 41580 800 41636 3388
rect 42028 3378 42084 3388
rect 42252 800 42308 4174
rect 43260 3666 43316 4620
rect 43708 4452 43764 4846
rect 44044 4452 44100 4462
rect 43708 4450 44100 4452
rect 43708 4398 44046 4450
rect 44098 4398 44100 4450
rect 43708 4396 44100 4398
rect 43260 3614 43262 3666
rect 43314 3614 43316 3666
rect 43260 3602 43316 3614
rect 44044 3220 44100 4396
rect 45388 4226 45444 6300
rect 45388 4174 45390 4226
rect 45442 4174 45444 4226
rect 45388 4162 45444 4174
rect 45948 4450 46004 4462
rect 45948 4398 45950 4450
rect 46002 4398 46004 4450
rect 45948 4228 46004 4398
rect 45948 4162 46004 4172
rect 46060 3668 46116 6636
rect 46172 5236 46228 5246
rect 46620 5236 46676 20076
rect 46172 5234 46676 5236
rect 46172 5182 46174 5234
rect 46226 5182 46676 5234
rect 46172 5180 46676 5182
rect 46172 5170 46228 5180
rect 46620 5122 46676 5180
rect 46620 5070 46622 5122
rect 46674 5070 46676 5122
rect 46620 5058 46676 5070
rect 46844 4564 46900 22204
rect 46956 22258 47012 22270
rect 46956 22206 46958 22258
rect 47010 22206 47012 22258
rect 46956 22036 47012 22206
rect 46956 21970 47012 21980
rect 47180 21700 47236 21710
rect 47180 21606 47236 21644
rect 46956 20132 47012 20142
rect 46956 20038 47012 20076
rect 47180 20020 47236 20030
rect 47180 19926 47236 19964
rect 47516 19796 47572 26012
rect 48076 24948 48132 27692
rect 48300 27188 48356 28476
rect 48300 27122 48356 27132
rect 47628 24946 48132 24948
rect 47628 24894 48078 24946
rect 48130 24894 48132 24946
rect 47628 24892 48132 24894
rect 47628 24722 47684 24892
rect 47628 24670 47630 24722
rect 47682 24670 47684 24722
rect 47628 24658 47684 24670
rect 47852 23716 47908 23726
rect 47852 23622 47908 23660
rect 47740 22260 47796 22270
rect 47740 22166 47796 22204
rect 47964 21812 48020 24892
rect 48076 24882 48132 24892
rect 48524 23716 48580 29150
rect 49420 29650 49476 31892
rect 49420 29598 49422 29650
rect 49474 29598 49476 29650
rect 49420 28532 49476 29598
rect 49420 28466 49476 28476
rect 49756 31892 50036 31948
rect 48524 23650 48580 23660
rect 48188 22484 48244 22494
rect 48188 22390 48244 22428
rect 48524 22484 48580 22494
rect 48524 22148 48580 22428
rect 48412 21812 48468 21822
rect 47964 21810 48468 21812
rect 47964 21758 48414 21810
rect 48466 21758 48468 21810
rect 47964 21756 48468 21758
rect 47964 21586 48020 21756
rect 47964 21534 47966 21586
rect 48018 21534 48020 21586
rect 47964 21522 48020 21534
rect 47628 20916 47684 20926
rect 47628 20822 47684 20860
rect 48300 20916 48356 21756
rect 48412 21746 48468 21756
rect 48300 20802 48356 20860
rect 48300 20750 48302 20802
rect 48354 20750 48356 20802
rect 48300 20738 48356 20750
rect 48524 20188 48580 22092
rect 48972 20916 49028 20926
rect 48972 20822 49028 20860
rect 48300 20132 48580 20188
rect 48300 20020 48356 20132
rect 48300 19926 48356 19964
rect 47516 19730 47572 19740
rect 47740 19906 47796 19918
rect 47740 19854 47742 19906
rect 47794 19854 47796 19906
rect 47740 19796 47796 19854
rect 47740 19730 47796 19740
rect 48076 5794 48132 5806
rect 48076 5742 48078 5794
rect 48130 5742 48132 5794
rect 47292 5236 47348 5246
rect 46284 4562 46900 4564
rect 46284 4510 46846 4562
rect 46898 4510 46900 4562
rect 46284 4508 46900 4510
rect 46284 4450 46340 4508
rect 46844 4498 46900 4508
rect 46956 5234 47348 5236
rect 46956 5182 47294 5234
rect 47346 5182 47348 5234
rect 46956 5180 47348 5182
rect 46284 4398 46286 4450
rect 46338 4398 46340 4450
rect 46284 4386 46340 4398
rect 46508 3668 46564 3678
rect 46060 3666 46564 3668
rect 46060 3614 46510 3666
rect 46562 3614 46564 3666
rect 46060 3612 46564 3614
rect 46508 3602 46564 3612
rect 44268 3444 44324 3454
rect 44268 3350 44324 3388
rect 45164 3444 45220 3454
rect 45388 3444 45444 3454
rect 45220 3442 45444 3444
rect 45220 3390 45390 3442
rect 45442 3390 45444 3442
rect 45220 3388 45444 3390
rect 43820 3164 44100 3220
rect 43820 800 43876 3164
rect 45164 800 45220 3388
rect 45388 3378 45444 3388
rect 46956 1428 47012 5180
rect 47292 5170 47348 5180
rect 48076 5012 48132 5742
rect 48524 5236 48580 5246
rect 48076 4946 48132 4956
rect 48412 5012 48468 5022
rect 48412 4918 48468 4956
rect 48524 4338 48580 5180
rect 49196 5236 49252 5246
rect 49196 5142 49252 5180
rect 49756 5236 49812 31892
rect 49756 5170 49812 5180
rect 50316 5234 50372 43484
rect 50428 43538 50484 43596
rect 50428 43486 50430 43538
rect 50482 43486 50484 43538
rect 50428 43474 50484 43486
rect 50764 43538 50820 43596
rect 50764 43486 50766 43538
rect 50818 43486 50820 43538
rect 50764 43474 50820 43486
rect 50428 43092 50484 43102
rect 50428 42866 50484 43036
rect 50428 42814 50430 42866
rect 50482 42814 50484 42866
rect 50428 42802 50484 42814
rect 50876 42866 50932 42878
rect 50876 42814 50878 42866
rect 50930 42814 50932 42866
rect 50540 42532 50596 42542
rect 50428 42530 50596 42532
rect 50428 42478 50542 42530
rect 50594 42478 50596 42530
rect 50428 42476 50596 42478
rect 50428 40628 50484 42476
rect 50540 42466 50596 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50876 41972 50932 42814
rect 50876 41906 50932 41916
rect 50988 41748 51044 44604
rect 51548 44548 51604 44558
rect 51324 44212 51380 44222
rect 51324 44118 51380 44156
rect 51548 42754 51604 44492
rect 51884 44322 51940 48972
rect 52108 48916 52164 48926
rect 52220 48916 52276 49196
rect 52108 48914 52388 48916
rect 52108 48862 52110 48914
rect 52162 48862 52388 48914
rect 52108 48860 52388 48862
rect 52108 48850 52164 48860
rect 51996 48804 52052 48814
rect 51996 48692 52052 48748
rect 51996 48636 52164 48692
rect 52108 48242 52164 48636
rect 52108 48190 52110 48242
rect 52162 48190 52164 48242
rect 52108 48178 52164 48190
rect 52220 46004 52276 46014
rect 52220 45668 52276 45948
rect 52220 45602 52276 45612
rect 52332 45332 52388 48860
rect 52444 48692 52500 48702
rect 52444 48242 52500 48636
rect 52444 48190 52446 48242
rect 52498 48190 52500 48242
rect 52444 46114 52500 48190
rect 52444 46062 52446 46114
rect 52498 46062 52500 46114
rect 52444 46050 52500 46062
rect 52444 45332 52500 45342
rect 52332 45330 52500 45332
rect 52332 45278 52446 45330
rect 52498 45278 52500 45330
rect 52332 45276 52500 45278
rect 52444 45266 52500 45276
rect 51996 45220 52052 45230
rect 51996 45126 52052 45164
rect 52556 44660 52612 51660
rect 52892 51490 52948 51884
rect 52892 51438 52894 51490
rect 52946 51438 52948 51490
rect 52892 51426 52948 51438
rect 52668 50708 52724 50718
rect 52668 50614 52724 50652
rect 53004 50428 53060 52444
rect 53116 51380 53172 54012
rect 53340 54012 53452 54068
rect 53228 52836 53284 52846
rect 53228 52742 53284 52780
rect 53340 52722 53396 54012
rect 53452 54002 53508 54012
rect 53564 53732 53620 56588
rect 53900 56420 53956 56430
rect 53788 56306 53844 56318
rect 53788 56254 53790 56306
rect 53842 56254 53844 56306
rect 53788 56084 53844 56254
rect 53788 56018 53844 56028
rect 53676 55972 53732 55982
rect 53676 55878 53732 55916
rect 53788 55858 53844 55870
rect 53788 55806 53790 55858
rect 53842 55806 53844 55858
rect 53788 55748 53844 55806
rect 53788 55682 53844 55692
rect 53900 55468 53956 56364
rect 53788 55412 53956 55468
rect 53676 55300 53732 55310
rect 53676 55206 53732 55244
rect 53788 54740 53844 55412
rect 53900 55298 53956 55310
rect 53900 55246 53902 55298
rect 53954 55246 53956 55298
rect 53900 55188 53956 55246
rect 53900 55122 53956 55132
rect 53900 54740 53956 54750
rect 53788 54738 53956 54740
rect 53788 54686 53902 54738
rect 53954 54686 53956 54738
rect 53788 54684 53956 54686
rect 53900 54674 53956 54684
rect 54012 53842 54068 56812
rect 54124 55412 54180 55422
rect 54124 55318 54180 55356
rect 54012 53790 54014 53842
rect 54066 53790 54068 53842
rect 54012 53778 54068 53790
rect 53564 53676 53956 53732
rect 53564 53396 53620 53406
rect 53340 52670 53342 52722
rect 53394 52670 53396 52722
rect 53340 52658 53396 52670
rect 53452 53284 53508 53294
rect 53340 51604 53396 51614
rect 53116 51378 53284 51380
rect 53116 51326 53118 51378
rect 53170 51326 53284 51378
rect 53116 51324 53284 51326
rect 53116 51314 53172 51324
rect 53004 50372 53172 50428
rect 52780 49700 52836 49710
rect 52668 49364 52724 49374
rect 52668 49138 52724 49308
rect 52668 49086 52670 49138
rect 52722 49086 52724 49138
rect 52668 49074 52724 49086
rect 52668 48916 52724 48926
rect 52668 47570 52724 48860
rect 52780 48244 52836 49644
rect 53004 48356 53060 48366
rect 53004 48262 53060 48300
rect 52780 48178 52836 48188
rect 52668 47518 52670 47570
rect 52722 47518 52724 47570
rect 52668 47506 52724 47518
rect 52668 46114 52724 46126
rect 52668 46062 52670 46114
rect 52722 46062 52724 46114
rect 52668 46004 52724 46062
rect 52668 46002 52948 46004
rect 52668 45950 52670 46002
rect 52722 45950 52948 46002
rect 52668 45948 52948 45950
rect 52668 45938 52724 45948
rect 52108 44604 52612 44660
rect 52108 44548 52164 44604
rect 51884 44270 51886 44322
rect 51938 44270 51940 44322
rect 51548 42702 51550 42754
rect 51602 42702 51604 42754
rect 51548 42644 51604 42702
rect 51772 44212 51828 44222
rect 51772 42756 51828 44156
rect 51772 42624 51828 42700
rect 51884 44100 51940 44270
rect 51884 43538 51940 44044
rect 51884 43486 51886 43538
rect 51938 43486 51940 43538
rect 51436 42532 51492 42542
rect 51436 42438 51492 42476
rect 50876 41692 51044 41748
rect 50540 41076 50596 41086
rect 50540 40982 50596 41020
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50428 40572 50708 40628
rect 50652 40290 50708 40572
rect 50652 40238 50654 40290
rect 50706 40238 50708 40290
rect 50652 40226 50708 40238
rect 50876 40626 50932 41692
rect 50876 40574 50878 40626
rect 50930 40574 50932 40626
rect 50876 40068 50932 40574
rect 50988 41076 51044 41086
rect 50988 40290 51044 41020
rect 51548 40626 51604 42588
rect 51884 41972 51940 43486
rect 51996 44546 52164 44548
rect 51996 44494 52110 44546
rect 52162 44494 52164 44546
rect 51996 44492 52164 44494
rect 51996 44436 52052 44492
rect 52108 44482 52164 44492
rect 51996 43426 52052 44380
rect 52444 44100 52500 44110
rect 52444 44006 52500 44044
rect 52892 43652 52948 45948
rect 53116 44212 53172 50372
rect 53228 50034 53284 51324
rect 53340 50818 53396 51548
rect 53340 50766 53342 50818
rect 53394 50766 53396 50818
rect 53340 50754 53396 50766
rect 53228 49982 53230 50034
rect 53282 49982 53284 50034
rect 53228 49364 53284 49982
rect 53228 49298 53284 49308
rect 53452 49138 53508 53228
rect 53564 51044 53620 53340
rect 53676 52948 53732 52958
rect 53676 52854 53732 52892
rect 53564 50978 53620 50988
rect 53676 52388 53732 52398
rect 53564 50818 53620 50830
rect 53564 50766 53566 50818
rect 53618 50766 53620 50818
rect 53564 50706 53620 50766
rect 53564 50654 53566 50706
rect 53618 50654 53620 50706
rect 53564 50642 53620 50654
rect 53676 50428 53732 52332
rect 53788 51938 53844 51950
rect 53788 51886 53790 51938
rect 53842 51886 53844 51938
rect 53788 50932 53844 51886
rect 53900 51828 53956 53676
rect 54012 53172 54068 53182
rect 54012 53058 54068 53116
rect 54012 53006 54014 53058
rect 54066 53006 54068 53058
rect 54012 52994 54068 53006
rect 53900 51762 53956 51772
rect 54012 52612 54068 52622
rect 53900 51604 53956 51614
rect 53900 51490 53956 51548
rect 53900 51438 53902 51490
rect 53954 51438 53956 51490
rect 53900 51426 53956 51438
rect 54012 51378 54068 52556
rect 54236 52052 54292 57820
rect 54572 57876 54628 58158
rect 54572 57810 54628 57820
rect 54348 57764 54404 57774
rect 54348 57670 54404 57708
rect 54684 57538 54740 57550
rect 54684 57486 54686 57538
rect 54738 57486 54740 57538
rect 54684 57428 54740 57486
rect 54684 57362 54740 57372
rect 54572 56754 54628 56766
rect 54572 56702 54574 56754
rect 54626 56702 54628 56754
rect 54460 56196 54516 56206
rect 54460 56102 54516 56140
rect 54572 55300 54628 56702
rect 55132 56532 55188 59388
rect 55468 59332 55524 59836
rect 55580 59332 55636 59342
rect 55468 59330 55636 59332
rect 55468 59278 55582 59330
rect 55634 59278 55636 59330
rect 55468 59276 55636 59278
rect 55580 59266 55636 59276
rect 54796 56476 55188 56532
rect 55244 59220 55300 59230
rect 55244 57538 55300 59164
rect 55244 57486 55246 57538
rect 55298 57486 55300 57538
rect 54684 55970 54740 55982
rect 54684 55918 54686 55970
rect 54738 55918 54740 55970
rect 54684 55636 54740 55918
rect 54684 55570 54740 55580
rect 54684 55300 54740 55310
rect 54572 55298 54740 55300
rect 54572 55246 54686 55298
rect 54738 55246 54740 55298
rect 54572 55244 54740 55246
rect 54684 55234 54740 55244
rect 54572 55074 54628 55086
rect 54572 55022 54574 55074
rect 54626 55022 54628 55074
rect 54572 54740 54628 55022
rect 54796 54964 54852 56476
rect 55020 56306 55076 56318
rect 55020 56254 55022 56306
rect 55074 56254 55076 56306
rect 54908 56084 54964 56094
rect 54908 55990 54964 56028
rect 55020 55522 55076 56254
rect 55020 55470 55022 55522
rect 55074 55470 55076 55522
rect 55020 55458 55076 55470
rect 55132 56082 55188 56094
rect 55132 56030 55134 56082
rect 55186 56030 55188 56082
rect 55132 55524 55188 56030
rect 55244 55748 55300 57486
rect 55356 58660 55412 58670
rect 55356 58324 55412 58604
rect 55580 58324 55636 58334
rect 55356 58322 55636 58324
rect 55356 58270 55582 58322
rect 55634 58270 55636 58322
rect 55356 58268 55636 58270
rect 55356 57540 55412 58268
rect 55580 58258 55636 58268
rect 55356 57474 55412 57484
rect 55468 57764 55524 57774
rect 55356 56420 55412 56430
rect 55356 56194 55412 56364
rect 55356 56142 55358 56194
rect 55410 56142 55412 56194
rect 55356 56130 55412 56142
rect 55244 55692 55412 55748
rect 55132 55458 55188 55468
rect 54908 55300 54964 55310
rect 55132 55300 55188 55310
rect 54908 55298 55188 55300
rect 54908 55246 54910 55298
rect 54962 55246 55134 55298
rect 55186 55246 55188 55298
rect 54908 55244 55188 55246
rect 54908 55234 54964 55244
rect 55132 55234 55188 55244
rect 55244 55074 55300 55086
rect 55244 55022 55246 55074
rect 55298 55022 55300 55074
rect 54796 54908 55188 54964
rect 54572 54684 55076 54740
rect 54572 54516 54628 54554
rect 54572 54450 54628 54460
rect 55020 54514 55076 54684
rect 55020 54462 55022 54514
rect 55074 54462 55076 54514
rect 55020 54450 55076 54462
rect 54348 54404 54404 54414
rect 54348 54310 54404 54348
rect 54572 54292 54628 54302
rect 54012 51326 54014 51378
rect 54066 51326 54068 51378
rect 54012 51314 54068 51326
rect 54124 52050 54292 52052
rect 54124 51998 54238 52050
rect 54290 51998 54292 52050
rect 54124 51996 54292 51998
rect 53788 50866 53844 50876
rect 53900 51268 53956 51278
rect 53900 50708 53956 51212
rect 54124 51156 54180 51996
rect 54236 51986 54292 51996
rect 54348 53060 54404 53070
rect 53452 49086 53454 49138
rect 53506 49086 53508 49138
rect 53452 49074 53508 49086
rect 53564 50372 53732 50428
rect 53788 50596 53844 50606
rect 53228 48132 53284 48142
rect 53228 45220 53284 48076
rect 53452 46562 53508 46574
rect 53452 46510 53454 46562
rect 53506 46510 53508 46562
rect 53452 46228 53508 46510
rect 53452 46162 53508 46172
rect 53228 45154 53284 45164
rect 53228 44996 53284 45006
rect 53228 44902 53284 44940
rect 53116 44146 53172 44156
rect 53564 44212 53620 50372
rect 53676 49924 53732 49934
rect 53676 49830 53732 49868
rect 53788 47570 53844 50540
rect 53900 49252 53956 50652
rect 54012 51100 54180 51156
rect 54012 49924 54068 51100
rect 54348 51044 54404 53004
rect 54460 52164 54516 52174
rect 54460 52070 54516 52108
rect 54012 49858 54068 49868
rect 54124 50988 54404 51044
rect 53900 49196 54068 49252
rect 53788 47518 53790 47570
rect 53842 47518 53844 47570
rect 53788 47506 53844 47518
rect 53900 49026 53956 49038
rect 53900 48974 53902 49026
rect 53954 48974 53956 49026
rect 53788 47234 53844 47246
rect 53788 47182 53790 47234
rect 53842 47182 53844 47234
rect 53676 46564 53732 46574
rect 53676 46002 53732 46508
rect 53676 45950 53678 46002
rect 53730 45950 53732 46002
rect 53676 45938 53732 45950
rect 53676 45220 53732 45230
rect 53676 45126 53732 45164
rect 53788 44996 53844 47182
rect 53900 46004 53956 48974
rect 54012 48916 54068 49196
rect 54124 49138 54180 50988
rect 54236 50818 54292 50830
rect 54236 50766 54238 50818
rect 54290 50766 54292 50818
rect 54236 50708 54292 50766
rect 54236 50642 54292 50652
rect 54572 50596 54628 54236
rect 54796 54292 54852 54302
rect 55132 54292 55188 54908
rect 54796 54290 55188 54292
rect 54796 54238 54798 54290
rect 54850 54238 55188 54290
rect 54796 54236 55188 54238
rect 54684 53284 54740 53294
rect 54684 53170 54740 53228
rect 54684 53118 54686 53170
rect 54738 53118 54740 53170
rect 54684 53106 54740 53118
rect 54796 53060 54852 54236
rect 54796 52994 54852 53004
rect 55244 52948 55300 55022
rect 55244 52882 55300 52892
rect 54796 52834 54852 52846
rect 54796 52782 54798 52834
rect 54850 52782 54852 52834
rect 54796 52388 54852 52782
rect 54796 52322 54852 52332
rect 54908 52722 54964 52734
rect 55356 52724 55412 55692
rect 55468 54516 55524 57708
rect 55580 57538 55636 57550
rect 55580 57486 55582 57538
rect 55634 57486 55636 57538
rect 55580 57204 55636 57486
rect 55580 57138 55636 57148
rect 55692 54516 55748 60508
rect 56028 60498 56084 60508
rect 55916 60004 55972 60014
rect 55916 60002 56084 60004
rect 55916 59950 55918 60002
rect 55970 59950 56084 60002
rect 55916 59948 56084 59950
rect 55916 59938 55972 59948
rect 55916 59220 55972 59230
rect 55916 59126 55972 59164
rect 55804 58996 55860 59006
rect 55804 58434 55860 58940
rect 56028 58546 56084 59948
rect 56028 58494 56030 58546
rect 56082 58494 56084 58546
rect 56028 58482 56084 58494
rect 55804 58382 55806 58434
rect 55858 58382 55860 58434
rect 55804 58370 55860 58382
rect 56028 58324 56084 58334
rect 56028 57874 56084 58268
rect 56028 57822 56030 57874
rect 56082 57822 56084 57874
rect 56028 57764 56084 57822
rect 56140 57876 56196 60732
rect 56476 60114 56532 61742
rect 56476 60062 56478 60114
rect 56530 60062 56532 60114
rect 56476 60050 56532 60062
rect 56252 59444 56308 59454
rect 56252 58434 56308 59388
rect 56364 59218 56420 59230
rect 56364 59166 56366 59218
rect 56418 59166 56420 59218
rect 56364 58772 56420 59166
rect 56364 58706 56420 58716
rect 56252 58382 56254 58434
rect 56306 58382 56308 58434
rect 56252 58370 56308 58382
rect 56588 58212 56644 63084
rect 56700 62468 56756 62478
rect 56700 62188 56756 62412
rect 56700 62132 56868 62188
rect 56812 61348 56868 62132
rect 56812 61346 56980 61348
rect 56812 61294 56814 61346
rect 56866 61294 56980 61346
rect 56812 61292 56980 61294
rect 56812 61282 56868 61292
rect 56924 60676 56980 61292
rect 56812 60004 56868 60014
rect 56700 59890 56756 59902
rect 56700 59838 56702 59890
rect 56754 59838 56756 59890
rect 56700 58324 56756 59838
rect 56812 58658 56868 59948
rect 56924 59892 56980 60620
rect 56924 59826 56980 59836
rect 57036 60002 57092 60014
rect 57036 59950 57038 60002
rect 57090 59950 57092 60002
rect 56812 58606 56814 58658
rect 56866 58606 56868 58658
rect 56812 58594 56868 58606
rect 56924 59668 56980 59678
rect 56924 58996 56980 59612
rect 57036 59444 57092 59950
rect 57148 59668 57204 64766
rect 57260 60228 57316 65548
rect 58492 65538 58548 65548
rect 57484 65380 57540 65390
rect 57372 65156 57428 65166
rect 57372 63250 57428 65100
rect 57484 64596 57540 65324
rect 57820 65380 57876 65390
rect 57820 64706 57876 65324
rect 58044 65378 58100 65390
rect 58044 65326 58046 65378
rect 58098 65326 58100 65378
rect 58044 65156 58100 65326
rect 58044 65090 58100 65100
rect 57820 64654 57822 64706
rect 57874 64654 57876 64706
rect 57820 64642 57876 64654
rect 57932 64820 57988 64830
rect 57484 64530 57540 64540
rect 57932 64594 57988 64764
rect 57932 64542 57934 64594
rect 57986 64542 57988 64594
rect 57932 64530 57988 64542
rect 57820 64148 57876 64158
rect 58380 64148 58436 64158
rect 58604 64148 58660 66444
rect 58940 66386 58996 66444
rect 58940 66334 58942 66386
rect 58994 66334 58996 66386
rect 58940 66322 58996 66334
rect 59052 67060 59108 67070
rect 58716 66276 58772 66286
rect 58716 65604 58772 66220
rect 58716 65538 58772 65548
rect 58828 64708 58884 64718
rect 58828 64614 58884 64652
rect 58940 64596 58996 64606
rect 58940 64502 58996 64540
rect 57596 63924 57652 63934
rect 57596 63830 57652 63868
rect 57372 63198 57374 63250
rect 57426 63198 57428 63250
rect 57372 63140 57428 63198
rect 57372 63074 57428 63084
rect 57708 63364 57764 63374
rect 57596 62242 57652 62254
rect 57596 62190 57598 62242
rect 57650 62190 57652 62242
rect 57596 62188 57652 62190
rect 57260 60162 57316 60172
rect 57484 62132 57652 62188
rect 57484 60004 57540 62132
rect 57484 59938 57540 59948
rect 57596 61348 57652 61358
rect 57708 61348 57764 63308
rect 57820 63250 57876 64092
rect 58268 64146 58660 64148
rect 58268 64094 58382 64146
rect 58434 64094 58660 64146
rect 58268 64092 58660 64094
rect 58268 63924 58324 64092
rect 58380 64082 58436 64092
rect 58268 63858 58324 63868
rect 58492 63924 58548 63934
rect 58492 63810 58548 63868
rect 59052 63922 59108 67004
rect 59052 63870 59054 63922
rect 59106 63870 59108 63922
rect 59052 63858 59108 63870
rect 58492 63758 58494 63810
rect 58546 63758 58548 63810
rect 58492 63746 58548 63758
rect 57820 63198 57822 63250
rect 57874 63198 57876 63250
rect 57820 63186 57876 63198
rect 58156 63698 58212 63710
rect 58156 63646 58158 63698
rect 58210 63646 58212 63698
rect 58156 62914 58212 63646
rect 58156 62862 58158 62914
rect 58210 62862 58212 62914
rect 58156 62850 58212 62862
rect 58268 63250 58324 63262
rect 58268 63198 58270 63250
rect 58322 63198 58324 63250
rect 58044 62468 58100 62478
rect 58044 62354 58100 62412
rect 58044 62302 58046 62354
rect 58098 62302 58100 62354
rect 58044 62290 58100 62302
rect 57596 61346 57764 61348
rect 57596 61294 57598 61346
rect 57650 61294 57764 61346
rect 57596 61292 57764 61294
rect 57820 61794 57876 61806
rect 57820 61742 57822 61794
rect 57874 61742 57876 61794
rect 57596 59892 57652 61292
rect 57820 61236 57876 61742
rect 58156 61460 58212 61470
rect 57708 61180 57876 61236
rect 58044 61346 58100 61358
rect 58044 61294 58046 61346
rect 58098 61294 58100 61346
rect 57708 60676 57764 61180
rect 58044 60900 58100 61294
rect 58044 60834 58100 60844
rect 57708 60582 57764 60620
rect 58156 60564 58212 61404
rect 57820 60004 57876 60014
rect 57820 59910 57876 59948
rect 57708 59892 57764 59902
rect 58156 59892 58212 60508
rect 58268 60340 58324 63198
rect 58940 63252 58996 63262
rect 58604 63140 58660 63150
rect 58940 63140 58996 63196
rect 58604 63046 58660 63084
rect 58828 63138 58996 63140
rect 58828 63086 58942 63138
rect 58994 63086 58996 63138
rect 58828 63084 58996 63086
rect 58492 63026 58548 63038
rect 58492 62974 58494 63026
rect 58546 62974 58548 63026
rect 58492 62466 58548 62974
rect 58492 62414 58494 62466
rect 58546 62414 58548 62466
rect 58492 62402 58548 62414
rect 58828 61794 58884 63084
rect 58940 63074 58996 63084
rect 59164 63140 59220 63150
rect 59164 63046 59220 63084
rect 58940 62468 58996 62478
rect 58940 62374 58996 62412
rect 58828 61742 58830 61794
rect 58882 61742 58884 61794
rect 58492 61348 58548 61358
rect 58492 61346 58772 61348
rect 58492 61294 58494 61346
rect 58546 61294 58772 61346
rect 58492 61292 58772 61294
rect 58492 61282 58548 61292
rect 58380 60900 58436 60910
rect 58380 60806 58436 60844
rect 58492 60788 58548 60798
rect 58492 60694 58548 60732
rect 58604 60564 58660 60574
rect 58604 60470 58660 60508
rect 58716 60452 58772 61292
rect 58828 60900 58884 61742
rect 59276 61682 59332 68236
rect 59388 66388 59444 102452
rect 59724 89572 59780 89582
rect 59724 89478 59780 89516
rect 60732 89572 60788 89582
rect 60732 73948 60788 89516
rect 59388 66256 59444 66332
rect 60508 73892 60788 73948
rect 60508 67620 60564 73892
rect 60620 67956 60676 67966
rect 60620 67862 60676 67900
rect 60508 66946 60564 67564
rect 60508 66894 60510 66946
rect 60562 66894 60564 66946
rect 60508 66500 60564 66894
rect 60508 65492 60564 66444
rect 60620 67060 60676 67070
rect 60620 66386 60676 67004
rect 60620 66334 60622 66386
rect 60674 66334 60676 66386
rect 60620 66322 60676 66334
rect 60172 65436 60564 65492
rect 59836 65378 59892 65390
rect 59836 65326 59838 65378
rect 59890 65326 59892 65378
rect 59836 64596 59892 65326
rect 60172 64820 60228 65436
rect 60172 64688 60228 64764
rect 60956 65380 61012 65390
rect 60620 64708 60676 64718
rect 60620 64614 60676 64652
rect 59724 64372 59780 64382
rect 59276 61630 59278 61682
rect 59330 61630 59332 61682
rect 58828 60834 58884 60844
rect 58940 61346 58996 61358
rect 58940 61294 58942 61346
rect 58994 61294 58996 61346
rect 58940 60564 58996 61294
rect 59276 61012 59332 61630
rect 59500 64260 59556 64270
rect 59500 61684 59556 64204
rect 59612 63140 59668 63150
rect 59612 63046 59668 63084
rect 59724 62242 59780 64316
rect 59836 64148 59892 64540
rect 59836 64082 59892 64092
rect 59836 63924 59892 63934
rect 59836 63830 59892 63868
rect 60956 63252 61012 65324
rect 60956 63186 61012 63196
rect 59724 62190 59726 62242
rect 59778 62190 59780 62242
rect 59724 62178 59780 62190
rect 60620 62468 60676 62478
rect 60284 61796 60340 61806
rect 59724 61684 59780 61694
rect 59556 61682 59780 61684
rect 59556 61630 59726 61682
rect 59778 61630 59780 61682
rect 59556 61628 59780 61630
rect 59500 61552 59556 61628
rect 59724 61618 59780 61628
rect 59388 61012 59444 61022
rect 60284 61012 60340 61740
rect 59276 61010 59444 61012
rect 59276 60958 59390 61010
rect 59442 60958 59444 61010
rect 59276 60956 59444 60958
rect 59388 60946 59444 60956
rect 59836 61010 60340 61012
rect 59836 60958 60286 61010
rect 60338 60958 60340 61010
rect 59836 60956 60340 60958
rect 59612 60900 59668 60910
rect 59612 60806 59668 60844
rect 59836 60898 59892 60956
rect 60284 60946 60340 60956
rect 59836 60846 59838 60898
rect 59890 60846 59892 60898
rect 59836 60834 59892 60846
rect 59164 60788 59220 60798
rect 59500 60788 59556 60798
rect 59220 60732 59444 60788
rect 59164 60694 59220 60732
rect 58940 60498 58996 60508
rect 59052 60676 59108 60686
rect 58268 60284 58660 60340
rect 58492 60114 58548 60126
rect 58492 60062 58494 60114
rect 58546 60062 58548 60114
rect 58492 60004 58548 60062
rect 58492 59938 58548 59948
rect 57596 59890 57764 59892
rect 57596 59838 57710 59890
rect 57762 59838 57764 59890
rect 57596 59836 57764 59838
rect 57708 59826 57764 59836
rect 57932 59836 58212 59892
rect 57148 59602 57204 59612
rect 57484 59778 57540 59790
rect 57484 59726 57486 59778
rect 57538 59726 57540 59778
rect 57484 59444 57540 59726
rect 57036 59378 57092 59388
rect 57148 59388 57540 59444
rect 57820 59444 57876 59454
rect 56924 58436 56980 58940
rect 56700 58258 56756 58268
rect 56812 58380 56980 58436
rect 56140 57810 56196 57820
rect 56364 58156 56644 58212
rect 56028 57698 56084 57708
rect 55916 56980 55972 56990
rect 55916 56084 55972 56924
rect 56140 56308 56196 56318
rect 56364 56308 56420 58156
rect 56700 57876 56756 57886
rect 56700 57782 56756 57820
rect 56700 56980 56756 56990
rect 56700 56886 56756 56924
rect 56700 56308 56756 56318
rect 56364 56252 56644 56308
rect 56140 56194 56196 56252
rect 56140 56142 56142 56194
rect 56194 56142 56196 56194
rect 56140 56130 56196 56142
rect 55468 54460 55636 54516
rect 55468 54290 55524 54302
rect 55468 54238 55470 54290
rect 55522 54238 55524 54290
rect 55468 53508 55524 54238
rect 55468 53442 55524 53452
rect 55580 53172 55636 54460
rect 55692 54450 55748 54460
rect 55804 56082 55972 56084
rect 55804 56030 55918 56082
rect 55970 56030 55972 56082
rect 55804 56028 55972 56030
rect 55804 55860 55860 56028
rect 55916 56018 55972 56028
rect 56476 56082 56532 56094
rect 56476 56030 56478 56082
rect 56530 56030 56532 56082
rect 56364 55972 56420 55982
rect 56364 55878 56420 55916
rect 54908 52670 54910 52722
rect 54962 52670 54964 52722
rect 54796 52162 54852 52174
rect 54796 52110 54798 52162
rect 54850 52110 54852 52162
rect 54796 50820 54852 52110
rect 54908 51828 54964 52670
rect 54908 51268 54964 51772
rect 54908 51202 54964 51212
rect 55132 52668 55412 52724
rect 55468 53170 55636 53172
rect 55468 53118 55582 53170
rect 55634 53118 55636 53170
rect 55468 53116 55636 53118
rect 54796 50754 54852 50764
rect 54572 50530 54628 50540
rect 54908 50708 54964 50718
rect 54908 50594 54964 50652
rect 54908 50542 54910 50594
rect 54962 50542 54964 50594
rect 54908 50530 54964 50542
rect 54348 50484 54404 50494
rect 54348 50482 54516 50484
rect 54348 50430 54350 50482
rect 54402 50430 54516 50482
rect 54348 50428 54516 50430
rect 54348 50418 54404 50428
rect 54236 50370 54292 50382
rect 54236 50318 54238 50370
rect 54290 50318 54292 50370
rect 54236 50036 54292 50318
rect 54460 50148 54516 50428
rect 54460 50036 54516 50092
rect 55020 50148 55076 50158
rect 54572 50036 54628 50046
rect 54460 50034 54628 50036
rect 54460 49982 54574 50034
rect 54626 49982 54628 50034
rect 54460 49980 54628 49982
rect 54236 49970 54292 49980
rect 54572 49970 54628 49980
rect 54348 49924 54404 49934
rect 54404 49868 54516 49924
rect 54236 49810 54292 49822
rect 54236 49758 54238 49810
rect 54290 49758 54292 49810
rect 54348 49792 54404 49868
rect 54236 49588 54292 49758
rect 54236 49522 54292 49532
rect 54124 49086 54126 49138
rect 54178 49086 54180 49138
rect 54124 49074 54180 49086
rect 54460 49140 54516 49868
rect 55020 49922 55076 50092
rect 55020 49870 55022 49922
rect 55074 49870 55076 49922
rect 55020 49858 55076 49870
rect 55132 49924 55188 52668
rect 55468 52388 55524 53116
rect 55580 53106 55636 53116
rect 55804 54402 55860 55804
rect 56028 55860 56084 55870
rect 55916 55074 55972 55086
rect 55916 55022 55918 55074
rect 55970 55022 55972 55074
rect 55916 54964 55972 55022
rect 55916 54898 55972 54908
rect 55804 54350 55806 54402
rect 55858 54350 55860 54402
rect 55356 52332 55524 52388
rect 55356 51492 55412 52332
rect 55468 52164 55524 52174
rect 55468 52162 55636 52164
rect 55468 52110 55470 52162
rect 55522 52110 55636 52162
rect 55468 52108 55636 52110
rect 55468 52098 55524 52108
rect 55244 51436 55356 51492
rect 55244 50482 55300 51436
rect 55356 51426 55412 51436
rect 55468 51716 55524 51726
rect 55468 51044 55524 51660
rect 55244 50430 55246 50482
rect 55298 50430 55300 50482
rect 55244 50418 55300 50430
rect 55356 50820 55412 50830
rect 55132 49858 55188 49868
rect 55244 50036 55300 50046
rect 54460 49074 54516 49084
rect 54684 49476 54740 49486
rect 54348 49028 54404 49038
rect 54236 48916 54292 48926
rect 54012 48914 54292 48916
rect 54012 48862 54238 48914
rect 54290 48862 54292 48914
rect 54012 48860 54292 48862
rect 54012 48132 54068 48142
rect 54012 47682 54068 48076
rect 54236 48132 54292 48860
rect 54236 48066 54292 48076
rect 54012 47630 54014 47682
rect 54066 47630 54068 47682
rect 54012 47618 54068 47630
rect 54348 46898 54404 48972
rect 54572 47684 54628 47694
rect 54572 47570 54628 47628
rect 54572 47518 54574 47570
rect 54626 47518 54628 47570
rect 54572 47506 54628 47518
rect 54348 46846 54350 46898
rect 54402 46846 54404 46898
rect 54348 46834 54404 46846
rect 54684 46788 54740 49420
rect 55244 49028 55300 49980
rect 55132 48914 55188 48926
rect 55132 48862 55134 48914
rect 55186 48862 55188 48914
rect 55244 48896 55300 48972
rect 55356 48914 55412 50764
rect 55468 50706 55524 50988
rect 55468 50654 55470 50706
rect 55522 50654 55524 50706
rect 55468 50642 55524 50654
rect 55580 50428 55636 52108
rect 55692 52162 55748 52174
rect 55692 52110 55694 52162
rect 55746 52110 55748 52162
rect 55692 51940 55748 52110
rect 55692 51874 55748 51884
rect 55468 50372 55636 50428
rect 55468 50036 55524 50372
rect 55468 49970 55524 49980
rect 55804 49812 55860 54350
rect 56028 52946 56084 55804
rect 56364 55300 56420 55310
rect 56252 55076 56308 55086
rect 56140 55074 56308 55076
rect 56140 55022 56254 55074
rect 56306 55022 56308 55074
rect 56140 55020 56308 55022
rect 56140 54290 56196 55020
rect 56252 55010 56308 55020
rect 56252 54404 56308 54414
rect 56364 54404 56420 55244
rect 56476 54516 56532 56030
rect 56476 54450 56532 54460
rect 56252 54402 56420 54404
rect 56252 54350 56254 54402
rect 56306 54350 56420 54402
rect 56252 54348 56420 54350
rect 56252 54338 56308 54348
rect 56140 54238 56142 54290
rect 56194 54238 56196 54290
rect 56140 54226 56196 54238
rect 56028 52894 56030 52946
rect 56082 52894 56084 52946
rect 56028 52882 56084 52894
rect 56252 53508 56308 53518
rect 56252 52946 56308 53452
rect 56252 52894 56254 52946
rect 56306 52894 56308 52946
rect 56252 52882 56308 52894
rect 56364 52724 56420 54348
rect 56252 52668 56420 52724
rect 56476 52722 56532 52734
rect 56476 52670 56478 52722
rect 56530 52670 56532 52722
rect 54796 48130 54852 48142
rect 54796 48078 54798 48130
rect 54850 48078 54852 48130
rect 54796 48020 54852 48078
rect 54796 47954 54852 47964
rect 55020 47682 55076 47694
rect 55020 47630 55022 47682
rect 55074 47630 55076 47682
rect 55020 47234 55076 47630
rect 55020 47182 55022 47234
rect 55074 47182 55076 47234
rect 54684 46732 54852 46788
rect 54684 46564 54740 46574
rect 54684 46470 54740 46508
rect 53900 45938 53956 45948
rect 54124 45892 54180 45902
rect 54124 45798 54180 45836
rect 54572 45890 54628 45902
rect 54572 45838 54574 45890
rect 54626 45838 54628 45890
rect 53788 44930 53844 44940
rect 54012 45332 54068 45342
rect 53676 44212 53732 44222
rect 53564 44210 53732 44212
rect 53564 44158 53678 44210
rect 53730 44158 53732 44210
rect 53564 44156 53732 44158
rect 53452 44100 53508 44110
rect 53452 44006 53508 44044
rect 53564 43708 53620 44156
rect 53676 44146 53732 44156
rect 53788 44210 53844 44222
rect 53788 44158 53790 44210
rect 53842 44158 53844 44210
rect 52892 43520 52948 43596
rect 53452 43652 53620 43708
rect 53788 43764 53844 44158
rect 53900 44212 53956 44222
rect 53900 44118 53956 44156
rect 53788 43698 53844 43708
rect 54012 43652 54068 45276
rect 54572 45332 54628 45838
rect 54572 45266 54628 45276
rect 54124 44994 54180 45006
rect 54124 44942 54126 44994
rect 54178 44942 54180 44994
rect 54124 44100 54180 44942
rect 54460 44994 54516 45006
rect 54460 44942 54462 44994
rect 54514 44942 54516 44994
rect 54236 44882 54292 44894
rect 54236 44830 54238 44882
rect 54290 44830 54292 44882
rect 54236 44434 54292 44830
rect 54460 44772 54516 44942
rect 54460 44706 54516 44716
rect 54572 44884 54628 44894
rect 54236 44382 54238 44434
rect 54290 44382 54292 44434
rect 54236 44370 54292 44382
rect 54124 44034 54180 44044
rect 54460 44212 54516 44222
rect 52444 43428 52500 43438
rect 51996 43374 51998 43426
rect 52050 43374 52052 43426
rect 51996 42196 52052 43374
rect 52108 43426 52500 43428
rect 52108 43374 52446 43426
rect 52498 43374 52500 43426
rect 52108 43372 52500 43374
rect 52108 42754 52164 43372
rect 52444 43362 52500 43372
rect 53452 43204 53508 43652
rect 53900 43596 54068 43652
rect 54236 43652 54292 43662
rect 53564 43540 53620 43550
rect 53900 43540 53956 43596
rect 54236 43558 54292 43596
rect 53564 43538 53956 43540
rect 53564 43486 53566 43538
rect 53618 43486 53956 43538
rect 53564 43484 53956 43486
rect 53564 43474 53620 43484
rect 52108 42702 52110 42754
rect 52162 42702 52164 42754
rect 52108 42690 52164 42702
rect 52220 42980 52276 42990
rect 52220 42866 52276 42924
rect 52220 42814 52222 42866
rect 52274 42814 52276 42866
rect 52220 42308 52276 42814
rect 53452 42868 53508 43148
rect 53452 42802 53508 42812
rect 52556 42754 52612 42766
rect 52556 42702 52558 42754
rect 52610 42702 52612 42754
rect 52220 42252 52388 42308
rect 51996 42140 52276 42196
rect 51884 41906 51940 41916
rect 51548 40574 51550 40626
rect 51602 40574 51604 40626
rect 51548 40516 51604 40574
rect 51548 40450 51604 40460
rect 52220 40404 52276 42140
rect 52332 40626 52388 42252
rect 52556 41748 52612 42702
rect 53452 42642 53508 42654
rect 53452 42590 53454 42642
rect 53506 42590 53508 42642
rect 52668 42532 52724 42542
rect 53452 42532 53508 42590
rect 53676 42644 53732 42654
rect 53676 42550 53732 42588
rect 53900 42644 53956 43484
rect 54236 42644 54292 42654
rect 53900 42642 54292 42644
rect 53900 42590 54238 42642
rect 54290 42590 54292 42642
rect 53900 42588 54292 42590
rect 52668 42530 53508 42532
rect 52668 42478 52670 42530
rect 52722 42478 53508 42530
rect 52668 42476 53508 42478
rect 53564 42530 53620 42542
rect 53564 42478 53566 42530
rect 53618 42478 53620 42530
rect 52668 42466 52724 42476
rect 52780 41860 52836 41870
rect 52780 41766 52836 41804
rect 53452 41860 53508 41870
rect 52556 41682 52612 41692
rect 52668 41298 52724 41310
rect 52668 41246 52670 41298
rect 52722 41246 52724 41298
rect 52668 41076 52724 41246
rect 53452 41188 53508 41804
rect 53564 41300 53620 42478
rect 53900 41860 53956 42588
rect 54236 42578 54292 42588
rect 54460 42420 54516 44156
rect 53900 41794 53956 41804
rect 54124 42364 54516 42420
rect 53564 41234 53620 41244
rect 52668 41010 52724 41020
rect 53116 41186 53508 41188
rect 53116 41134 53454 41186
rect 53506 41134 53508 41186
rect 53116 41132 53508 41134
rect 52332 40574 52334 40626
rect 52386 40574 52388 40626
rect 52332 40562 52388 40574
rect 53116 40626 53172 41132
rect 53116 40574 53118 40626
rect 53170 40574 53172 40626
rect 53116 40562 53172 40574
rect 52668 40404 52724 40414
rect 52220 40402 52724 40404
rect 52220 40350 52670 40402
rect 52722 40350 52724 40402
rect 52220 40348 52724 40350
rect 52668 40338 52724 40348
rect 50988 40238 50990 40290
rect 51042 40238 51044 40290
rect 50988 40226 51044 40238
rect 50876 40012 51380 40068
rect 51324 39730 51380 40012
rect 51324 39678 51326 39730
rect 51378 39678 51380 39730
rect 51324 39666 51380 39678
rect 53340 39730 53396 41132
rect 53452 41122 53508 41132
rect 53564 41076 53620 41086
rect 53564 40068 53620 41020
rect 54124 40626 54180 42364
rect 54572 42196 54628 44828
rect 54796 44548 54852 46732
rect 55020 46564 55076 47182
rect 55132 46788 55188 48862
rect 55356 48862 55358 48914
rect 55410 48862 55412 48914
rect 55244 48244 55300 48254
rect 55244 48150 55300 48188
rect 55356 47682 55412 48862
rect 55356 47630 55358 47682
rect 55410 47630 55412 47682
rect 55356 47618 55412 47630
rect 55468 49756 55860 49812
rect 55916 52388 55972 52398
rect 55132 46732 55300 46788
rect 55020 46498 55076 46508
rect 55132 46562 55188 46574
rect 55132 46510 55134 46562
rect 55186 46510 55188 46562
rect 55132 46452 55188 46510
rect 54908 45332 54964 45342
rect 55132 45332 55188 46396
rect 54908 45330 55188 45332
rect 54908 45278 54910 45330
rect 54962 45278 55188 45330
rect 54908 45276 55188 45278
rect 54908 45266 54964 45276
rect 54348 42140 54628 42196
rect 54684 44492 54852 44548
rect 55020 44882 55076 44894
rect 55020 44830 55022 44882
rect 55074 44830 55076 44882
rect 54236 41300 54292 41310
rect 54236 41206 54292 41244
rect 54124 40574 54126 40626
rect 54178 40574 54180 40626
rect 54124 40562 54180 40574
rect 53676 40516 53732 40526
rect 53676 40422 53732 40460
rect 53564 40012 53732 40068
rect 53340 39678 53342 39730
rect 53394 39678 53396 39730
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 52780 38164 52836 38174
rect 53340 38164 53396 39678
rect 52780 38162 53396 38164
rect 52780 38110 52782 38162
rect 52834 38110 53396 38162
rect 52780 38108 53396 38110
rect 52780 38098 52836 38108
rect 53340 38052 53396 38108
rect 53564 38834 53620 38846
rect 53564 38782 53566 38834
rect 53618 38782 53620 38834
rect 53452 38052 53508 38062
rect 53340 38050 53508 38052
rect 53340 37998 53454 38050
rect 53506 37998 53508 38050
rect 53340 37996 53508 37998
rect 53452 37986 53508 37996
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 53564 37492 53620 38782
rect 53564 37426 53620 37436
rect 53564 37154 53620 37166
rect 53564 37102 53566 37154
rect 53618 37102 53620 37154
rect 53564 37044 53620 37102
rect 53564 36978 53620 36988
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 53676 15204 53732 40012
rect 53788 38946 53844 38958
rect 53788 38894 53790 38946
rect 53842 38894 53844 38946
rect 53788 38668 53844 38894
rect 53788 38612 54292 38668
rect 54236 38162 54292 38612
rect 54236 38110 54238 38162
rect 54290 38110 54292 38162
rect 54236 38098 54292 38110
rect 54236 37492 54292 37502
rect 54236 37398 54292 37436
rect 54348 26908 54404 42140
rect 54460 41860 54516 41870
rect 54460 40626 54516 41804
rect 54460 40574 54462 40626
rect 54514 40574 54516 40626
rect 54460 40562 54516 40574
rect 54684 38668 54740 44492
rect 55020 44322 55076 44830
rect 55244 44772 55300 46732
rect 55356 46004 55412 46014
rect 55356 45910 55412 45948
rect 55356 45668 55412 45678
rect 55356 44994 55412 45612
rect 55468 45220 55524 49756
rect 55916 48916 55972 52332
rect 56252 52052 56308 52668
rect 56364 52388 56420 52398
rect 56476 52388 56532 52670
rect 56364 52386 56532 52388
rect 56364 52334 56366 52386
rect 56418 52334 56532 52386
rect 56364 52332 56532 52334
rect 56364 52322 56420 52332
rect 56252 51986 56308 51996
rect 56364 51940 56420 51950
rect 56364 51602 56420 51884
rect 56364 51550 56366 51602
rect 56418 51550 56420 51602
rect 56364 51538 56420 51550
rect 56476 51828 56532 51838
rect 56140 51492 56196 51502
rect 56140 50594 56196 51436
rect 56140 50542 56142 50594
rect 56194 50542 56196 50594
rect 56140 50530 56196 50542
rect 56252 51490 56308 51502
rect 56252 51438 56254 51490
rect 56306 51438 56308 51490
rect 56252 49700 56308 51438
rect 56476 51490 56532 51772
rect 56476 51438 56478 51490
rect 56530 51438 56532 51490
rect 56476 51426 56532 51438
rect 56476 50932 56532 50942
rect 56476 50706 56532 50876
rect 56476 50654 56478 50706
rect 56530 50654 56532 50706
rect 56476 50642 56532 50654
rect 56252 49634 56308 49644
rect 56364 49924 56420 49934
rect 56364 49810 56420 49868
rect 56364 49758 56366 49810
rect 56418 49758 56420 49810
rect 55916 48860 56308 48916
rect 55804 48804 55860 48814
rect 55804 48802 56084 48804
rect 55804 48750 55806 48802
rect 55858 48750 56084 48802
rect 55804 48748 56084 48750
rect 55804 48738 55860 48748
rect 55692 48130 55748 48142
rect 55692 48078 55694 48130
rect 55746 48078 55748 48130
rect 55580 47460 55636 47470
rect 55692 47460 55748 48078
rect 56028 47682 56084 48748
rect 56140 48132 56196 48170
rect 56140 48066 56196 48076
rect 56028 47630 56030 47682
rect 56082 47630 56084 47682
rect 56028 47618 56084 47630
rect 56140 47908 56196 47918
rect 55580 47458 55748 47460
rect 55580 47406 55582 47458
rect 55634 47406 55748 47458
rect 55580 47404 55748 47406
rect 55916 47460 55972 47470
rect 55580 47394 55636 47404
rect 55804 46786 55860 46798
rect 55804 46734 55806 46786
rect 55858 46734 55860 46786
rect 55692 46450 55748 46462
rect 55692 46398 55694 46450
rect 55746 46398 55748 46450
rect 55692 46004 55748 46398
rect 55692 45938 55748 45948
rect 55804 45220 55860 46734
rect 55916 46452 55972 47404
rect 56028 47234 56084 47246
rect 56028 47182 56030 47234
rect 56082 47182 56084 47234
rect 56028 46786 56084 47182
rect 56028 46734 56030 46786
rect 56082 46734 56084 46786
rect 56028 46722 56084 46734
rect 55916 46386 55972 46396
rect 55468 45164 55636 45220
rect 55356 44942 55358 44994
rect 55410 44942 55412 44994
rect 55356 44884 55412 44942
rect 55356 44818 55412 44828
rect 55468 44996 55524 45006
rect 55244 44706 55300 44716
rect 55020 44270 55022 44322
rect 55074 44270 55076 44322
rect 55020 44258 55076 44270
rect 54796 44210 54852 44222
rect 54796 44158 54798 44210
rect 54850 44158 54852 44210
rect 54796 44100 54852 44158
rect 55356 44210 55412 44222
rect 55356 44158 55358 44210
rect 55410 44158 55412 44210
rect 54796 44034 54852 44044
rect 55132 44098 55188 44110
rect 55132 44046 55134 44098
rect 55186 44046 55188 44098
rect 55132 43652 55188 44046
rect 55356 43988 55412 44158
rect 55356 43922 55412 43932
rect 55132 43586 55188 43596
rect 55244 43876 55300 43886
rect 54908 43428 54964 43438
rect 54908 42868 54964 43372
rect 54908 42774 54964 42812
rect 54796 41972 54852 41982
rect 55244 41972 55300 43820
rect 55356 43764 55412 43774
rect 55356 42866 55412 43708
rect 55356 42814 55358 42866
rect 55410 42814 55412 42866
rect 55356 42802 55412 42814
rect 54796 41970 55300 41972
rect 54796 41918 54798 41970
rect 54850 41918 55246 41970
rect 55298 41918 55300 41970
rect 54796 41916 55300 41918
rect 54796 41906 54852 41916
rect 55244 41906 55300 41916
rect 54684 38612 54852 38668
rect 54572 37268 54628 37278
rect 54572 37174 54628 37212
rect 53676 15110 53732 15148
rect 54012 26852 54404 26908
rect 54684 37156 54740 37166
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50316 5182 50318 5234
rect 50370 5182 50372 5234
rect 48748 4900 48804 4910
rect 48748 4898 48916 4900
rect 48748 4846 48750 4898
rect 48802 4846 48916 4898
rect 48748 4844 48916 4846
rect 48748 4834 48804 4844
rect 48524 4286 48526 4338
rect 48578 4286 48580 4338
rect 48524 4274 48580 4286
rect 47404 4228 47460 4238
rect 46844 1372 47012 1428
rect 47180 4226 47460 4228
rect 47180 4174 47406 4226
rect 47458 4174 47460 4226
rect 47180 4172 47460 4174
rect 46508 812 46676 868
rect 46508 800 46564 812
rect 41580 728 41832 800
rect 42252 728 42504 800
rect 40264 200 40488 728
rect 41608 200 41832 728
rect 42280 200 42504 728
rect 43624 728 43876 800
rect 44968 728 45220 800
rect 46312 728 46564 800
rect 46620 756 46676 812
rect 46844 756 46900 1372
rect 47180 800 47236 4172
rect 47404 4162 47460 4172
rect 48524 3668 48580 3678
rect 48524 800 48580 3612
rect 48860 3554 48916 4844
rect 49420 4564 49476 4574
rect 49420 4470 49476 4508
rect 50316 4564 50372 5182
rect 54012 5012 54068 26852
rect 54460 15428 54516 15438
rect 54460 15334 54516 15372
rect 54124 15314 54180 15326
rect 54124 15262 54126 15314
rect 54178 15262 54180 15314
rect 54124 15204 54180 15262
rect 54124 15138 54180 15148
rect 54012 4946 54068 4956
rect 54460 4898 54516 4910
rect 54460 4846 54462 4898
rect 54514 4846 54516 4898
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 51660 4564 51716 4574
rect 50372 4508 50708 4564
rect 49980 4452 50036 4462
rect 49868 4450 50036 4452
rect 49868 4398 49982 4450
rect 50034 4398 50036 4450
rect 50316 4432 50372 4508
rect 50652 4450 50708 4508
rect 49868 4396 50036 4398
rect 49532 3668 49588 3678
rect 49532 3574 49588 3612
rect 48860 3502 48862 3554
rect 48914 3502 48916 3554
rect 48860 3490 48916 3502
rect 49868 800 49924 4396
rect 49980 4386 50036 4396
rect 50652 4398 50654 4450
rect 50706 4398 50708 4450
rect 50652 4386 50708 4398
rect 50988 4450 51044 4462
rect 50988 4398 50990 4450
rect 51042 4398 51044 4450
rect 50988 4340 51044 4398
rect 51548 4340 51604 4350
rect 50988 4338 51604 4340
rect 50988 4286 51550 4338
rect 51602 4286 51604 4338
rect 50988 4284 51604 4286
rect 51548 4274 51604 4284
rect 51660 3554 51716 4508
rect 53452 4450 53508 4462
rect 53452 4398 53454 4450
rect 53506 4398 53508 4450
rect 52220 4228 52276 4238
rect 51660 3502 51662 3554
rect 51714 3502 51716 3554
rect 51660 3490 51716 3502
rect 51884 4226 52276 4228
rect 51884 4174 52222 4226
rect 52274 4174 52276 4226
rect 51884 4172 52276 4174
rect 50764 3444 50820 3454
rect 50428 3442 50820 3444
rect 50428 3390 50766 3442
rect 50818 3390 50820 3442
rect 50428 3388 50820 3390
rect 50428 800 50484 3388
rect 50764 3378 50820 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51884 800 51940 4172
rect 52220 4162 52276 4172
rect 53116 3444 53172 3454
rect 53452 3444 53508 4398
rect 54460 4116 54516 4846
rect 54460 4050 54516 4060
rect 54572 4228 54628 4238
rect 53116 3442 53508 3444
rect 53116 3390 53118 3442
rect 53170 3390 53508 3442
rect 53116 3388 53508 3390
rect 53116 800 53172 3388
rect 54572 800 54628 4172
rect 54684 4226 54740 37100
rect 54796 20188 54852 38612
rect 55132 37828 55188 37838
rect 54908 37378 54964 37390
rect 54908 37326 54910 37378
rect 54962 37326 54964 37378
rect 54908 37044 54964 37326
rect 55132 37378 55188 37772
rect 55132 37326 55134 37378
rect 55186 37326 55188 37378
rect 55132 37314 55188 37326
rect 55468 37156 55524 44940
rect 55580 40292 55636 45164
rect 55804 45154 55860 45164
rect 55916 44996 55972 45006
rect 55916 44902 55972 44940
rect 55692 44772 55748 44782
rect 55692 42644 55748 44716
rect 56140 44548 56196 47852
rect 56252 47570 56308 48860
rect 56364 48804 56420 49758
rect 56476 49028 56532 49038
rect 56476 48934 56532 48972
rect 56364 48738 56420 48748
rect 56252 47518 56254 47570
rect 56306 47518 56308 47570
rect 56252 47506 56308 47518
rect 56364 47684 56420 47694
rect 56364 46900 56420 47628
rect 56476 47348 56532 47358
rect 56588 47348 56644 56252
rect 56700 54740 56756 56252
rect 56812 55410 56868 58380
rect 56812 55358 56814 55410
rect 56866 55358 56868 55410
rect 56812 55346 56868 55358
rect 56924 58210 56980 58222
rect 56924 58158 56926 58210
rect 56978 58158 56980 58210
rect 56700 54608 56756 54684
rect 56924 54516 56980 58158
rect 57036 58210 57092 58222
rect 57036 58158 57038 58210
rect 57090 58158 57092 58210
rect 57036 57764 57092 58158
rect 57036 57698 57092 57708
rect 56924 54450 56980 54460
rect 57036 57540 57092 57550
rect 56924 54292 56980 54302
rect 57036 54292 57092 57484
rect 56924 54290 57092 54292
rect 56924 54238 56926 54290
rect 56978 54238 57092 54290
rect 56924 54236 57092 54238
rect 56924 53172 56980 54236
rect 56700 52946 56756 52958
rect 56700 52894 56702 52946
rect 56754 52894 56756 52946
rect 56700 52724 56756 52894
rect 56700 52658 56756 52668
rect 56812 52948 56868 52958
rect 56812 52274 56868 52892
rect 56812 52222 56814 52274
rect 56866 52222 56868 52274
rect 56812 52210 56868 52222
rect 56700 51492 56756 51502
rect 56700 48466 56756 51436
rect 56924 51268 56980 53116
rect 56924 51202 56980 51212
rect 57036 52052 57092 52062
rect 56812 50372 56868 50382
rect 56812 49810 56868 50316
rect 56812 49758 56814 49810
rect 56866 49758 56868 49810
rect 56812 49588 56868 49758
rect 56812 49522 56868 49532
rect 56924 48804 56980 48814
rect 56924 48710 56980 48748
rect 56700 48414 56702 48466
rect 56754 48414 56756 48466
rect 56700 47684 56756 48414
rect 56700 47618 56756 47628
rect 56812 48132 56868 48142
rect 56476 47346 56756 47348
rect 56476 47294 56478 47346
rect 56530 47294 56756 47346
rect 56476 47292 56756 47294
rect 56476 47282 56532 47292
rect 56588 46900 56644 46910
rect 56364 46898 56644 46900
rect 56364 46846 56590 46898
rect 56642 46846 56644 46898
rect 56364 46844 56644 46846
rect 56588 46834 56644 46844
rect 56588 46452 56644 46462
rect 56364 45332 56420 45342
rect 56364 45238 56420 45276
rect 55916 44492 56196 44548
rect 55916 44434 55972 44492
rect 55916 44382 55918 44434
rect 55970 44382 55972 44434
rect 55916 44370 55972 44382
rect 55804 43988 55860 43998
rect 55804 42868 55860 43932
rect 56364 43428 56420 43438
rect 56364 43334 56420 43372
rect 55916 42868 55972 42878
rect 55804 42866 55972 42868
rect 55804 42814 55918 42866
rect 55970 42814 55972 42866
rect 55804 42812 55972 42814
rect 55916 42802 55972 42812
rect 56364 42868 56420 42878
rect 56588 42868 56644 46396
rect 56700 44434 56756 47292
rect 56812 45330 56868 48076
rect 57036 48132 57092 51996
rect 57036 48066 57092 48076
rect 56812 45278 56814 45330
rect 56866 45278 56868 45330
rect 56812 45266 56868 45278
rect 56700 44382 56702 44434
rect 56754 44382 56756 44434
rect 56700 44370 56756 44382
rect 57148 45108 57204 59388
rect 57820 59350 57876 59388
rect 57596 59332 57652 59342
rect 57596 59330 57764 59332
rect 57596 59278 57598 59330
rect 57650 59278 57764 59330
rect 57596 59276 57764 59278
rect 57596 59266 57652 59276
rect 57484 59218 57540 59230
rect 57484 59166 57486 59218
rect 57538 59166 57540 59218
rect 57484 58772 57540 59166
rect 57484 58706 57540 58716
rect 57596 58996 57652 59006
rect 57596 58436 57652 58940
rect 57484 58380 57652 58436
rect 57372 57764 57428 57774
rect 57372 57428 57428 57708
rect 57484 57650 57540 58380
rect 57484 57598 57486 57650
rect 57538 57598 57540 57650
rect 57484 57586 57540 57598
rect 57596 57762 57652 57774
rect 57596 57710 57598 57762
rect 57650 57710 57652 57762
rect 57372 57372 57540 57428
rect 57260 56980 57316 56990
rect 57260 56866 57316 56924
rect 57260 56814 57262 56866
rect 57314 56814 57316 56866
rect 57260 56802 57316 56814
rect 57372 56642 57428 56654
rect 57372 56590 57374 56642
rect 57426 56590 57428 56642
rect 57372 56308 57428 56590
rect 57372 56242 57428 56252
rect 57484 55410 57540 57372
rect 57596 56866 57652 57710
rect 57596 56814 57598 56866
rect 57650 56814 57652 56866
rect 57596 56802 57652 56814
rect 57708 56308 57764 59276
rect 57932 58436 57988 59836
rect 58492 59780 58548 59790
rect 58492 59686 58548 59724
rect 58156 59668 58212 59678
rect 58044 58436 58100 58446
rect 57932 58434 58100 58436
rect 57932 58382 58046 58434
rect 58098 58382 58100 58434
rect 57932 58380 58100 58382
rect 57820 58322 57876 58334
rect 57820 58270 57822 58322
rect 57874 58270 57876 58322
rect 57820 57652 57876 58270
rect 57820 57204 57876 57596
rect 57820 57138 57876 57148
rect 57932 56644 57988 58380
rect 58044 58370 58100 58380
rect 58044 56980 58100 56990
rect 58156 56980 58212 59612
rect 58492 59444 58548 59454
rect 58492 59330 58548 59388
rect 58492 59278 58494 59330
rect 58546 59278 58548 59330
rect 58492 59266 58548 59278
rect 58604 58660 58660 60284
rect 58716 60226 58772 60396
rect 58716 60174 58718 60226
rect 58770 60174 58772 60226
rect 58716 60162 58772 60174
rect 59052 59332 59108 60620
rect 59388 60228 59444 60732
rect 59500 60694 59556 60732
rect 59500 60228 59556 60238
rect 59388 60226 59556 60228
rect 59388 60174 59502 60226
rect 59554 60174 59556 60226
rect 59388 60172 59556 60174
rect 59500 60162 59556 60172
rect 59948 60228 60004 60238
rect 59948 60134 60004 60172
rect 59388 60004 59444 60042
rect 59388 59938 59444 59948
rect 59724 60004 59780 60014
rect 59724 59910 59780 59948
rect 60508 60004 60564 60014
rect 59388 59780 59444 59790
rect 60060 59780 60116 59790
rect 59388 59778 59556 59780
rect 59388 59726 59390 59778
rect 59442 59726 59556 59778
rect 59388 59724 59556 59726
rect 59388 59714 59444 59724
rect 58828 59330 59108 59332
rect 58828 59278 59054 59330
rect 59106 59278 59108 59330
rect 58828 59276 59108 59278
rect 58604 58594 58660 58604
rect 58716 59218 58772 59230
rect 58716 59166 58718 59218
rect 58770 59166 58772 59218
rect 58716 59108 58772 59166
rect 58268 58436 58324 58446
rect 58268 58342 58324 58380
rect 58380 58322 58436 58334
rect 58380 58270 58382 58322
rect 58434 58270 58436 58322
rect 58380 58212 58436 58270
rect 58380 57428 58436 58156
rect 58380 57362 58436 57372
rect 58716 58324 58772 59052
rect 58044 56978 58156 56980
rect 58044 56926 58046 56978
rect 58098 56926 58156 56978
rect 58044 56924 58156 56926
rect 58044 56914 58100 56924
rect 58156 56848 58212 56924
rect 58492 56980 58548 56990
rect 58716 56980 58772 58268
rect 58492 56978 58772 56980
rect 58492 56926 58494 56978
rect 58546 56926 58772 56978
rect 58492 56924 58772 56926
rect 58492 56914 58548 56924
rect 57932 56588 58660 56644
rect 57932 56308 57988 56318
rect 57708 56306 57988 56308
rect 57708 56254 57934 56306
rect 57986 56254 57988 56306
rect 57708 56252 57988 56254
rect 57596 56084 57652 56094
rect 57596 55990 57652 56028
rect 57484 55358 57486 55410
rect 57538 55358 57540 55410
rect 57484 55346 57540 55358
rect 57484 55076 57540 55086
rect 57372 52836 57428 52846
rect 57372 52742 57428 52780
rect 57484 52612 57540 55020
rect 57596 54516 57652 54526
rect 57596 54422 57652 54460
rect 57708 53172 57764 56252
rect 57932 56242 57988 56252
rect 58604 56306 58660 56588
rect 58604 56254 58606 56306
rect 58658 56254 58660 56306
rect 58604 56242 58660 56254
rect 57932 55298 57988 55310
rect 57932 55246 57934 55298
rect 57986 55246 57988 55298
rect 57932 55076 57988 55246
rect 58268 55186 58324 55198
rect 58828 55188 58884 59276
rect 59052 59266 59108 59276
rect 58940 59106 58996 59118
rect 58940 59054 58942 59106
rect 58994 59054 58996 59106
rect 58940 58434 58996 59054
rect 59276 58772 59332 58782
rect 58940 58382 58942 58434
rect 58994 58382 58996 58434
rect 58940 58370 58996 58382
rect 59164 58436 59220 58446
rect 59164 58342 59220 58380
rect 59052 58210 59108 58222
rect 59052 58158 59054 58210
rect 59106 58158 59108 58210
rect 58940 56980 58996 56990
rect 58940 56886 58996 56924
rect 59052 56194 59108 58158
rect 59276 57652 59332 58716
rect 59388 58660 59444 58670
rect 59388 58566 59444 58604
rect 59500 57876 59556 59724
rect 59948 59444 60004 59454
rect 59724 59442 60004 59444
rect 59724 59390 59950 59442
rect 60002 59390 60004 59442
rect 59724 59388 60004 59390
rect 59612 59218 59668 59230
rect 59612 59166 59614 59218
rect 59666 59166 59668 59218
rect 59612 58884 59668 59166
rect 59612 58818 59668 58828
rect 59612 58660 59668 58670
rect 59724 58660 59780 59388
rect 59948 59378 60004 59388
rect 59948 59220 60004 59230
rect 60060 59220 60116 59724
rect 60508 59778 60564 59948
rect 60508 59726 60510 59778
rect 60562 59726 60564 59778
rect 60508 59556 60564 59726
rect 60508 59490 60564 59500
rect 59948 59218 60116 59220
rect 59948 59166 59950 59218
rect 60002 59166 60116 59218
rect 59948 59164 60116 59166
rect 60284 59220 60340 59230
rect 60284 59218 60452 59220
rect 60284 59166 60286 59218
rect 60338 59166 60452 59218
rect 60284 59164 60452 59166
rect 59948 59154 60004 59164
rect 60284 59154 60340 59164
rect 59612 58658 59780 58660
rect 59612 58606 59614 58658
rect 59666 58606 59780 58658
rect 59612 58604 59780 58606
rect 59948 58660 60004 58670
rect 59612 58594 59668 58604
rect 59500 57820 59780 57876
rect 59276 56980 59332 57596
rect 59500 57650 59556 57662
rect 59500 57598 59502 57650
rect 59554 57598 59556 57650
rect 59500 57540 59556 57598
rect 59500 57474 59556 57484
rect 59276 56848 59332 56924
rect 59052 56142 59054 56194
rect 59106 56142 59108 56194
rect 59052 56130 59108 56142
rect 59724 56194 59780 57820
rect 59724 56142 59726 56194
rect 59778 56142 59780 56194
rect 59724 56130 59780 56142
rect 59836 56980 59892 56990
rect 59276 56082 59332 56094
rect 59276 56030 59278 56082
rect 59330 56030 59332 56082
rect 59164 55860 59220 55870
rect 59164 55766 59220 55804
rect 58268 55134 58270 55186
rect 58322 55134 58324 55186
rect 57932 55010 57988 55020
rect 58156 55076 58212 55086
rect 58156 54982 58212 55020
rect 58268 54964 58324 55134
rect 58716 55132 58884 55188
rect 58940 55636 58996 55646
rect 58940 55410 58996 55580
rect 58940 55358 58942 55410
rect 58994 55358 58996 55410
rect 58268 54898 58324 54908
rect 58604 55076 58660 55086
rect 57820 54740 57876 54750
rect 57820 54514 57876 54684
rect 57820 54462 57822 54514
rect 57874 54462 57876 54514
rect 57820 54292 57876 54462
rect 57820 54226 57876 54236
rect 58044 54516 58100 54526
rect 57932 53844 57988 53854
rect 57708 53106 57764 53116
rect 57820 53620 57876 53630
rect 57708 52836 57764 52846
rect 57708 52742 57764 52780
rect 57484 52556 57764 52612
rect 57260 52388 57316 52398
rect 57260 52274 57316 52332
rect 57260 52222 57262 52274
rect 57314 52222 57316 52274
rect 57260 52210 57316 52222
rect 57708 52274 57764 52556
rect 57708 52222 57710 52274
rect 57762 52222 57764 52274
rect 57708 52210 57764 52222
rect 57484 51492 57540 51502
rect 57484 51398 57540 51436
rect 57708 51492 57764 51502
rect 57708 51378 57764 51436
rect 57708 51326 57710 51378
rect 57762 51326 57764 51378
rect 57708 51314 57764 51326
rect 57708 50820 57764 50830
rect 57484 49028 57540 49066
rect 57372 48972 57484 49028
rect 57260 48244 57316 48254
rect 57260 45668 57316 48188
rect 57372 47682 57428 48972
rect 57484 48962 57540 48972
rect 57708 49026 57764 50764
rect 57708 48974 57710 49026
rect 57762 48974 57764 49026
rect 57372 47630 57374 47682
rect 57426 47630 57428 47682
rect 57372 47618 57428 47630
rect 57484 48804 57540 48814
rect 57372 47460 57428 47470
rect 57372 47366 57428 47404
rect 57372 46900 57428 46910
rect 57484 46900 57540 48748
rect 57596 48244 57652 48254
rect 57596 48150 57652 48188
rect 57708 47908 57764 48974
rect 57596 47852 57764 47908
rect 57820 49810 57876 53564
rect 57932 53170 57988 53788
rect 57932 53118 57934 53170
rect 57986 53118 57988 53170
rect 57932 53106 57988 53118
rect 58044 53058 58100 54460
rect 58492 54516 58548 54526
rect 58492 54422 58548 54460
rect 58492 53508 58548 53518
rect 58492 53396 58548 53452
rect 58268 53340 58548 53396
rect 58044 53006 58046 53058
rect 58098 53006 58100 53058
rect 58044 52994 58100 53006
rect 58156 53284 58212 53294
rect 58156 52946 58212 53228
rect 58156 52894 58158 52946
rect 58210 52894 58212 52946
rect 57820 49758 57822 49810
rect 57874 49758 57876 49810
rect 57596 47012 57652 47852
rect 57708 47682 57764 47694
rect 57708 47630 57710 47682
rect 57762 47630 57764 47682
rect 57708 47570 57764 47630
rect 57708 47518 57710 47570
rect 57762 47518 57764 47570
rect 57708 47348 57764 47518
rect 57708 47282 57764 47292
rect 57596 46946 57652 46956
rect 57372 46898 57540 46900
rect 57372 46846 57374 46898
rect 57426 46846 57540 46898
rect 57372 46844 57540 46846
rect 57372 46834 57428 46844
rect 57260 45602 57316 45612
rect 57484 46564 57540 46574
rect 57484 45330 57540 46508
rect 57596 45668 57652 45678
rect 57596 45574 57652 45612
rect 57484 45278 57486 45330
rect 57538 45278 57540 45330
rect 57484 45266 57540 45278
rect 57820 45332 57876 49758
rect 57932 52612 57988 52622
rect 57932 45892 57988 52556
rect 58044 52500 58100 52510
rect 58156 52500 58212 52894
rect 58100 52444 58212 52500
rect 58044 51602 58100 52444
rect 58156 52276 58212 52286
rect 58268 52276 58324 53340
rect 58156 52274 58324 52276
rect 58156 52222 58158 52274
rect 58210 52222 58324 52274
rect 58156 52220 58324 52222
rect 58156 52210 58212 52220
rect 58044 51550 58046 51602
rect 58098 51550 58100 51602
rect 58044 51538 58100 51550
rect 58268 51380 58324 52220
rect 58380 53172 58436 53182
rect 58380 52500 58436 53116
rect 58492 53170 58548 53340
rect 58492 53118 58494 53170
rect 58546 53118 58548 53170
rect 58492 53106 58548 53118
rect 58604 52612 58660 55020
rect 58716 54180 58772 55132
rect 58828 54964 58884 54974
rect 58828 54292 58884 54908
rect 58940 54852 58996 55358
rect 59164 55300 59220 55310
rect 59164 55206 59220 55244
rect 59052 55076 59108 55086
rect 59276 55076 59332 56030
rect 59500 56084 59556 56094
rect 59556 56028 59668 56084
rect 59500 55952 59556 56028
rect 59388 55412 59444 55422
rect 59388 55318 59444 55356
rect 59052 55074 59332 55076
rect 59052 55022 59054 55074
rect 59106 55022 59332 55074
rect 59052 55020 59332 55022
rect 59500 55298 59556 55310
rect 59500 55246 59502 55298
rect 59554 55246 59556 55298
rect 59500 55076 59556 55246
rect 59052 55010 59108 55020
rect 59500 55010 59556 55020
rect 59612 54852 59668 56028
rect 59836 55412 59892 56924
rect 59948 56978 60004 58604
rect 60396 58210 60452 59164
rect 60396 58158 60398 58210
rect 60450 58158 60452 58210
rect 59948 56926 59950 56978
rect 60002 56926 60004 56978
rect 59948 56914 60004 56926
rect 60172 57538 60228 57550
rect 60172 57486 60174 57538
rect 60226 57486 60228 57538
rect 60060 56644 60116 56654
rect 60060 56550 60116 56588
rect 60172 56306 60228 57486
rect 60396 56868 60452 58158
rect 60620 57764 60676 62412
rect 60732 60676 60788 60686
rect 60732 60674 60900 60676
rect 60732 60622 60734 60674
rect 60786 60622 60900 60674
rect 60732 60620 60900 60622
rect 60732 60610 60788 60620
rect 60620 57632 60676 57708
rect 60844 60564 60900 60620
rect 60844 58994 60900 60508
rect 60956 60228 61012 60238
rect 60956 59442 61012 60172
rect 60956 59390 60958 59442
rect 61010 59390 61012 59442
rect 60956 59378 61012 59390
rect 60844 58942 60846 58994
rect 60898 58942 60900 58994
rect 60396 56802 60452 56812
rect 60508 57540 60564 57550
rect 60172 56254 60174 56306
rect 60226 56254 60228 56306
rect 60172 56084 60228 56254
rect 60172 55748 60228 56028
rect 60172 55682 60228 55692
rect 60060 55412 60116 55422
rect 59836 55410 60116 55412
rect 59836 55358 60062 55410
rect 60114 55358 60116 55410
rect 59836 55356 60116 55358
rect 60060 55346 60116 55356
rect 58940 54796 59220 54852
rect 59164 54738 59220 54796
rect 59164 54686 59166 54738
rect 59218 54686 59220 54738
rect 59164 54674 59220 54686
rect 59276 54796 59668 54852
rect 59276 54516 59332 54796
rect 59164 54460 59332 54516
rect 59388 54684 60116 54740
rect 59388 54514 59444 54684
rect 59388 54462 59390 54514
rect 59442 54462 59444 54514
rect 59052 54292 59108 54302
rect 58828 54290 59108 54292
rect 58828 54238 59054 54290
rect 59106 54238 59108 54290
rect 58828 54236 59108 54238
rect 59052 54180 59108 54236
rect 58716 54124 58884 54180
rect 58716 53730 58772 53742
rect 58716 53678 58718 53730
rect 58770 53678 58772 53730
rect 58716 53620 58772 53678
rect 58716 53554 58772 53564
rect 58828 53172 58884 54124
rect 59052 54114 59108 54124
rect 58716 52948 58772 52958
rect 58716 52854 58772 52892
rect 58604 52546 58660 52556
rect 58380 51716 58436 52444
rect 58828 52388 58884 53116
rect 59164 52612 59220 54460
rect 59388 54450 59444 54462
rect 59948 54514 60004 54526
rect 59948 54462 59950 54514
rect 60002 54462 60004 54514
rect 59836 54180 59892 54190
rect 59612 53956 59668 53966
rect 59612 53862 59668 53900
rect 59276 53844 59332 53854
rect 59276 53750 59332 53788
rect 59836 53844 59892 54124
rect 59724 53732 59780 53742
rect 59500 53506 59556 53518
rect 59500 53454 59502 53506
rect 59554 53454 59556 53506
rect 59388 53172 59444 53182
rect 59388 53078 59444 53116
rect 59500 53060 59556 53454
rect 59500 52994 59556 53004
rect 59276 52836 59332 52846
rect 59276 52742 59332 52780
rect 59612 52724 59668 52734
rect 59500 52722 59668 52724
rect 59500 52670 59614 52722
rect 59666 52670 59668 52722
rect 59500 52668 59668 52670
rect 59164 52556 59332 52612
rect 58828 52322 58884 52332
rect 58828 51940 58884 51950
rect 58828 51846 58884 51884
rect 58940 51938 58996 51950
rect 58940 51886 58942 51938
rect 58994 51886 58996 51938
rect 58940 51828 58996 51886
rect 58940 51762 58996 51772
rect 59052 51938 59108 51950
rect 59052 51886 59054 51938
rect 59106 51886 59108 51938
rect 58380 51660 58884 51716
rect 58828 51602 58884 51660
rect 58828 51550 58830 51602
rect 58882 51550 58884 51602
rect 58604 51492 58660 51502
rect 58604 51398 58660 51436
rect 58268 51324 58436 51380
rect 58380 50372 58436 51324
rect 58492 50820 58548 50830
rect 58492 50706 58548 50764
rect 58492 50654 58494 50706
rect 58546 50654 58548 50706
rect 58492 50642 58548 50654
rect 58828 50708 58884 51550
rect 58380 50306 58436 50316
rect 58604 50594 58660 50606
rect 58828 50596 58884 50652
rect 58604 50542 58606 50594
rect 58658 50542 58660 50594
rect 58044 48802 58100 48814
rect 58044 48750 58046 48802
rect 58098 48750 58100 48802
rect 58044 47908 58100 48750
rect 58604 48804 58660 50542
rect 58716 50540 58884 50596
rect 58940 51378 58996 51390
rect 58940 51326 58942 51378
rect 58994 51326 58996 51378
rect 58716 49028 58772 50540
rect 58828 50372 58884 50382
rect 58828 49476 58884 50316
rect 58828 49138 58884 49420
rect 58828 49086 58830 49138
rect 58882 49086 58884 49138
rect 58828 49074 58884 49086
rect 58716 48962 58772 48972
rect 58940 48916 58996 51326
rect 59052 49700 59108 51886
rect 59052 49634 59108 49644
rect 59164 51940 59220 51950
rect 59164 50932 59220 51884
rect 59164 49364 59220 50876
rect 59276 50428 59332 52556
rect 59388 52052 59444 52062
rect 59388 51958 59444 51996
rect 59388 51604 59444 51614
rect 59500 51604 59556 52668
rect 59612 52658 59668 52668
rect 59388 51602 59556 51604
rect 59388 51550 59390 51602
rect 59442 51550 59556 51602
rect 59388 51548 59556 51550
rect 59388 51538 59444 51548
rect 59388 50708 59444 50718
rect 59388 50614 59444 50652
rect 59500 50484 59556 51548
rect 59724 51604 59780 53676
rect 59724 51538 59780 51548
rect 59724 50596 59780 50606
rect 59836 50596 59892 53788
rect 59948 51380 60004 54462
rect 60060 53508 60116 54684
rect 60508 53844 60564 57484
rect 60844 57540 60900 58942
rect 60844 57474 60900 57484
rect 60732 56644 60788 56654
rect 60732 56550 60788 56588
rect 61068 56308 61124 116508
rect 61740 116338 61796 116508
rect 61740 116286 61742 116338
rect 61794 116286 61796 116338
rect 61740 116274 61796 116286
rect 62636 115780 62692 119200
rect 63980 117010 64036 119200
rect 63980 116958 63982 117010
rect 64034 116958 64036 117010
rect 63980 116946 64036 116958
rect 65212 117010 65268 117022
rect 65212 116958 65214 117010
rect 65266 116958 65268 117010
rect 65212 116562 65268 116958
rect 65212 116510 65214 116562
rect 65266 116510 65268 116562
rect 65212 116498 65268 116510
rect 65324 116564 65380 119200
rect 67228 117010 67284 117022
rect 67228 116958 67230 117010
rect 67282 116958 67284 117010
rect 65916 116844 66180 116854
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 65916 116778 66180 116788
rect 65324 116498 65380 116508
rect 66444 116564 66500 116574
rect 66444 116470 66500 116508
rect 64540 116452 64596 116462
rect 63868 116450 64596 116452
rect 63868 116398 64542 116450
rect 64594 116398 64596 116450
rect 63868 116396 64596 116398
rect 62860 115780 62916 115790
rect 62636 115778 62916 115780
rect 62636 115726 62862 115778
rect 62914 115726 62916 115778
rect 62636 115724 62916 115726
rect 62860 115714 62916 115724
rect 62972 115780 63028 115790
rect 62972 114994 63028 115724
rect 62972 114942 62974 114994
rect 63026 114942 63028 114994
rect 62972 114884 63028 114942
rect 62972 114818 63028 114828
rect 63644 114882 63700 114894
rect 63644 114830 63646 114882
rect 63698 114830 63700 114882
rect 61292 114660 61348 114670
rect 61292 94388 61348 114604
rect 63644 114324 63700 114830
rect 63868 114770 63924 116396
rect 64540 116386 64596 116396
rect 67228 115890 67284 116958
rect 67340 116564 67396 119200
rect 68684 117572 68740 119200
rect 68684 117516 68852 117572
rect 67340 116498 67396 116508
rect 68460 117010 68516 117022
rect 68460 116958 68462 117010
rect 68514 116958 68516 117010
rect 67564 116452 67620 116462
rect 67564 116450 68404 116452
rect 67564 116398 67566 116450
rect 67618 116398 68404 116450
rect 67564 116396 68404 116398
rect 67564 116386 67620 116396
rect 68348 116116 68404 116396
rect 68460 116450 68516 116958
rect 68460 116398 68462 116450
rect 68514 116398 68516 116450
rect 68460 116386 68516 116398
rect 68348 116060 68740 116116
rect 67228 115838 67230 115890
rect 67282 115838 67284 115890
rect 67228 115826 67284 115838
rect 68684 115890 68740 116060
rect 68684 115838 68686 115890
rect 68738 115838 68740 115890
rect 68684 115826 68740 115838
rect 68796 115892 68852 117516
rect 69132 116564 69188 116574
rect 69132 116470 69188 116508
rect 70588 116562 70644 119200
rect 70588 116510 70590 116562
rect 70642 116510 70644 116562
rect 70588 116498 70644 116510
rect 71372 116452 71428 116462
rect 71260 116450 71428 116452
rect 71260 116398 71374 116450
rect 71426 116398 71428 116450
rect 71260 116396 71428 116398
rect 68796 115826 68852 115836
rect 69580 115892 69636 115902
rect 69580 115798 69636 115836
rect 63980 115666 64036 115678
rect 63980 115614 63982 115666
rect 64034 115614 64036 115666
rect 63980 115556 64036 115614
rect 67004 115666 67060 115678
rect 67004 115614 67006 115666
rect 67058 115614 67060 115666
rect 64428 115556 64484 115566
rect 63980 115554 64484 115556
rect 63980 115502 64430 115554
rect 64482 115502 64484 115554
rect 63980 115500 64484 115502
rect 63868 114718 63870 114770
rect 63922 114718 63924 114770
rect 63868 114706 63924 114718
rect 63644 114258 63700 114268
rect 64092 114324 64148 114362
rect 64092 114258 64148 114268
rect 61292 94322 61348 94332
rect 61852 93604 61908 93614
rect 61852 73948 61908 93548
rect 61628 73892 61908 73948
rect 61964 86436 62020 86446
rect 61964 73948 62020 86380
rect 62188 77812 62244 77822
rect 61964 73892 62132 73948
rect 61404 67956 61460 67966
rect 61292 67060 61348 67070
rect 61292 66966 61348 67004
rect 61180 64036 61236 64046
rect 61180 61684 61236 63980
rect 61404 63252 61460 67900
rect 61628 67956 61684 73892
rect 61628 67844 61684 67900
rect 61852 67844 61908 67854
rect 61628 67842 61908 67844
rect 61628 67790 61854 67842
rect 61906 67790 61908 67842
rect 61628 67788 61908 67790
rect 61852 67778 61908 67788
rect 61516 67618 61572 67630
rect 62076 67620 62132 73892
rect 62188 68180 62244 77756
rect 63084 68516 63140 68526
rect 62188 68114 62244 68124
rect 62636 68514 63140 68516
rect 62636 68462 63086 68514
rect 63138 68462 63140 68514
rect 62636 68460 63140 68462
rect 62636 67842 62692 68460
rect 63084 68450 63140 68460
rect 63980 68514 64036 68526
rect 63980 68462 63982 68514
rect 64034 68462 64036 68514
rect 62636 67790 62638 67842
rect 62690 67790 62692 67842
rect 62524 67732 62580 67742
rect 62524 67638 62580 67676
rect 61516 67566 61518 67618
rect 61570 67566 61572 67618
rect 61516 66274 61572 67566
rect 61516 66222 61518 66274
rect 61570 66222 61572 66274
rect 61516 66210 61572 66222
rect 61628 67564 62132 67620
rect 61516 65492 61572 65502
rect 61516 65398 61572 65436
rect 61404 63196 61572 63252
rect 61404 63028 61460 63038
rect 61404 62934 61460 62972
rect 61516 62804 61572 63196
rect 61180 61618 61236 61628
rect 61404 62748 61572 62804
rect 61292 60788 61348 60798
rect 61292 60694 61348 60732
rect 61292 60228 61348 60238
rect 61292 60114 61348 60172
rect 61292 60062 61294 60114
rect 61346 60062 61348 60114
rect 61292 60050 61348 60062
rect 61180 59220 61236 59258
rect 61180 59154 61236 59164
rect 61404 58436 61460 62748
rect 61516 62356 61572 62366
rect 61516 61010 61572 62300
rect 61516 60958 61518 61010
rect 61570 60958 61572 61010
rect 61516 60946 61572 60958
rect 61404 58100 61460 58380
rect 61404 58034 61460 58044
rect 61516 59668 61572 59678
rect 61404 56980 61460 56990
rect 61404 56644 61460 56924
rect 61516 56868 61572 59612
rect 61628 59332 61684 67564
rect 62076 67060 62132 67070
rect 61964 66948 62020 66958
rect 61740 66946 62020 66948
rect 61740 66894 61966 66946
rect 62018 66894 62020 66946
rect 61740 66892 62020 66894
rect 61740 66162 61796 66892
rect 61964 66882 62020 66892
rect 61740 66110 61742 66162
rect 61794 66110 61796 66162
rect 61740 66098 61796 66110
rect 62076 65604 62132 67004
rect 62636 66724 62692 67790
rect 63644 67954 63700 67966
rect 63644 67902 63646 67954
rect 63698 67902 63700 67954
rect 63308 67730 63364 67742
rect 63308 67678 63310 67730
rect 63362 67678 63364 67730
rect 62188 66050 62244 66062
rect 62188 65998 62190 66050
rect 62242 65998 62244 66050
rect 62188 65828 62244 65998
rect 62188 65772 62580 65828
rect 62300 65604 62356 65614
rect 62076 65548 62244 65604
rect 62188 64930 62244 65548
rect 62300 65510 62356 65548
rect 62412 65492 62468 65502
rect 62412 65398 62468 65436
rect 62524 65490 62580 65772
rect 62524 65438 62526 65490
rect 62578 65438 62580 65490
rect 62524 65268 62580 65438
rect 62188 64878 62190 64930
rect 62242 64878 62244 64930
rect 62188 64818 62244 64878
rect 62188 64766 62190 64818
rect 62242 64766 62244 64818
rect 62188 64754 62244 64766
rect 62412 65212 62580 65268
rect 61964 64036 62020 64046
rect 61964 63810 62020 63980
rect 61964 63758 61966 63810
rect 62018 63758 62020 63810
rect 61964 63746 62020 63758
rect 62412 63252 62468 65212
rect 62636 65156 62692 66668
rect 62972 67060 63028 67070
rect 62972 66274 63028 67004
rect 62972 66222 62974 66274
rect 63026 66222 63028 66274
rect 62972 66210 63028 66222
rect 63308 65714 63364 67678
rect 63532 67618 63588 67630
rect 63532 67566 63534 67618
rect 63586 67566 63588 67618
rect 63532 67172 63588 67566
rect 63532 67106 63588 67116
rect 63644 66388 63700 67902
rect 63980 67172 64036 68462
rect 63756 66388 63812 66398
rect 63644 66386 63812 66388
rect 63644 66334 63758 66386
rect 63810 66334 63812 66386
rect 63644 66332 63812 66334
rect 63756 66322 63812 66332
rect 63308 65662 63310 65714
rect 63362 65662 63364 65714
rect 63308 65650 63364 65662
rect 63532 65940 63588 65950
rect 62972 65492 63028 65502
rect 62972 65490 63140 65492
rect 62972 65438 62974 65490
rect 63026 65438 63140 65490
rect 62972 65436 63140 65438
rect 62972 65426 63028 65436
rect 62636 65100 63028 65156
rect 62076 63196 62468 63252
rect 62524 64930 62580 64942
rect 62524 64878 62526 64930
rect 62578 64878 62580 64930
rect 62076 63028 62132 63196
rect 61852 62916 61908 62926
rect 61852 62914 62020 62916
rect 61852 62862 61854 62914
rect 61906 62862 62020 62914
rect 61852 62860 62020 62862
rect 61852 62850 61908 62860
rect 61852 62356 61908 62394
rect 61852 62290 61908 62300
rect 61964 62188 62020 62860
rect 62076 62804 62132 62972
rect 62188 63028 62244 63038
rect 62412 63028 62468 63038
rect 62188 63026 62468 63028
rect 62188 62974 62190 63026
rect 62242 62974 62414 63026
rect 62466 62974 62468 63026
rect 62188 62972 62468 62974
rect 62188 62962 62244 62972
rect 62412 62962 62468 62972
rect 62076 62748 62356 62804
rect 61740 62132 62020 62188
rect 61740 60898 61796 62132
rect 61740 60846 61742 60898
rect 61794 60846 61796 60898
rect 61740 60834 61796 60846
rect 61852 60900 61908 60910
rect 61852 60114 61908 60844
rect 61964 60788 62020 60798
rect 61964 60694 62020 60732
rect 61852 60062 61854 60114
rect 61906 60062 61908 60114
rect 61852 59444 61908 60062
rect 62300 60226 62356 62748
rect 62524 62580 62580 64878
rect 62636 64820 62692 64830
rect 62636 64036 62692 64764
rect 62860 64484 62916 64494
rect 62748 64036 62804 64046
rect 62692 64034 62804 64036
rect 62692 63982 62750 64034
rect 62802 63982 62804 64034
rect 62692 63980 62804 63982
rect 62636 63904 62692 63980
rect 62748 63970 62804 63980
rect 62860 63476 62916 64428
rect 62524 62354 62580 62524
rect 62524 62302 62526 62354
rect 62578 62302 62580 62354
rect 62524 61682 62580 62302
rect 62524 61630 62526 61682
rect 62578 61630 62580 61682
rect 62524 61618 62580 61630
rect 62636 63420 62916 63476
rect 62412 60788 62468 60798
rect 62412 60694 62468 60732
rect 62300 60174 62302 60226
rect 62354 60174 62356 60226
rect 62300 60114 62356 60174
rect 62300 60062 62302 60114
rect 62354 60062 62356 60114
rect 62300 60050 62356 60062
rect 61852 59378 61908 59388
rect 62636 59556 62692 63420
rect 62860 63250 62916 63262
rect 62860 63198 62862 63250
rect 62914 63198 62916 63250
rect 62748 63028 62804 63038
rect 62860 63028 62916 63198
rect 62972 63140 63028 65100
rect 63084 65044 63140 65436
rect 63196 65380 63252 65390
rect 63196 65286 63252 65324
rect 63532 65378 63588 65884
rect 63980 65604 64036 67116
rect 64092 67956 64148 67966
rect 64204 67956 64260 115500
rect 64428 115490 64484 115500
rect 64764 115556 64820 115566
rect 64428 114884 64484 114894
rect 64428 114790 64484 114828
rect 64764 114770 64820 115500
rect 64764 114718 64766 114770
rect 64818 114718 64820 114770
rect 64764 114706 64820 114718
rect 65212 115556 65268 115566
rect 64092 67954 64260 67956
rect 64092 67902 64094 67954
rect 64146 67902 64260 67954
rect 64092 67900 64260 67902
rect 65212 114324 65268 115500
rect 66332 115556 66388 115566
rect 66332 115462 66388 115500
rect 67004 115556 67060 115614
rect 65916 115276 66180 115286
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 65916 115210 66180 115220
rect 67004 114996 67060 115500
rect 69020 115666 69076 115678
rect 69020 115614 69022 115666
rect 69074 115614 69076 115666
rect 69020 115444 69076 115614
rect 70700 115668 70756 115678
rect 70140 115554 70196 115566
rect 70140 115502 70142 115554
rect 70194 115502 70196 115554
rect 69020 115378 69076 115388
rect 69580 115444 69636 115454
rect 67004 114930 67060 114940
rect 64092 67732 64148 67900
rect 64092 66946 64148 67676
rect 64540 67618 64596 67630
rect 64540 67566 64542 67618
rect 64594 67566 64596 67618
rect 64540 67172 64596 67566
rect 64540 67106 64596 67116
rect 64092 66894 64094 66946
rect 64146 66894 64148 66946
rect 64092 66882 64148 66894
rect 64540 66946 64596 66958
rect 64540 66894 64542 66946
rect 64594 66894 64596 66946
rect 63980 65538 64036 65548
rect 64092 66052 64148 66062
rect 63532 65326 63534 65378
rect 63586 65326 63588 65378
rect 63532 65314 63588 65326
rect 63868 65380 63924 65390
rect 63084 64988 63476 65044
rect 63420 64818 63476 64988
rect 63420 64766 63422 64818
rect 63474 64766 63476 64818
rect 63420 64754 63476 64766
rect 63644 64706 63700 64718
rect 63644 64654 63646 64706
rect 63698 64654 63700 64706
rect 63084 64260 63140 64270
rect 63084 64146 63140 64204
rect 63084 64094 63086 64146
rect 63138 64094 63140 64146
rect 63084 64082 63140 64094
rect 63644 63812 63700 64654
rect 63868 64484 63924 65324
rect 64092 64706 64148 65996
rect 64540 65940 64596 66894
rect 64540 65874 64596 65884
rect 64652 66052 64708 66062
rect 64652 65490 64708 65996
rect 64652 65438 64654 65490
rect 64706 65438 64708 65490
rect 64652 65426 64708 65438
rect 64988 65604 65044 65614
rect 64092 64654 64094 64706
rect 64146 64654 64148 64706
rect 64092 64642 64148 64654
rect 63868 64418 63924 64428
rect 64092 64372 64148 64382
rect 63868 64148 63924 64158
rect 63196 63810 63700 63812
rect 63196 63758 63646 63810
rect 63698 63758 63700 63810
rect 63196 63756 63700 63758
rect 63196 63362 63252 63756
rect 63644 63746 63700 63756
rect 63756 63812 63812 63822
rect 63756 63718 63812 63756
rect 63196 63310 63198 63362
rect 63250 63310 63252 63362
rect 63196 63298 63252 63310
rect 62972 63084 63252 63140
rect 62748 63026 62916 63028
rect 62748 62974 62750 63026
rect 62802 62974 62916 63026
rect 62748 62972 62916 62974
rect 62748 62962 62804 62972
rect 62972 62916 63028 62926
rect 62972 62822 63028 62860
rect 63084 62580 63140 62590
rect 63084 61684 63140 62524
rect 63196 62188 63252 63084
rect 63756 62916 63812 62926
rect 63756 62578 63812 62860
rect 63868 62914 63924 64092
rect 63980 63698 64036 63710
rect 63980 63646 63982 63698
rect 64034 63646 64036 63698
rect 63980 63588 64036 63646
rect 63980 63522 64036 63532
rect 63868 62862 63870 62914
rect 63922 62862 63924 62914
rect 63868 62850 63924 62862
rect 63756 62526 63758 62578
rect 63810 62526 63812 62578
rect 63756 62514 63812 62526
rect 64092 62580 64148 64316
rect 64876 64036 64932 64046
rect 64204 63924 64260 63934
rect 64204 63028 64260 63868
rect 64764 63922 64820 63934
rect 64764 63870 64766 63922
rect 64818 63870 64820 63922
rect 64764 63812 64820 63870
rect 64316 63028 64372 63038
rect 64204 63026 64372 63028
rect 64204 62974 64318 63026
rect 64370 62974 64372 63026
rect 64204 62972 64372 62974
rect 64316 62962 64372 62972
rect 64764 62916 64820 63756
rect 64764 62850 64820 62860
rect 64652 62580 64708 62590
rect 64092 62578 64708 62580
rect 64092 62526 64654 62578
rect 64706 62526 64708 62578
rect 64092 62524 64708 62526
rect 63644 62356 63700 62366
rect 63700 62300 63812 62356
rect 63644 62262 63700 62300
rect 63196 62132 63476 62188
rect 63084 61628 63252 61684
rect 62972 60674 63028 60686
rect 62972 60622 62974 60674
rect 63026 60622 63028 60674
rect 62972 59890 63028 60622
rect 62972 59838 62974 59890
rect 63026 59838 63028 59890
rect 62972 59826 63028 59838
rect 63084 60226 63140 60238
rect 63084 60174 63086 60226
rect 63138 60174 63140 60226
rect 62860 59778 62916 59790
rect 62860 59726 62862 59778
rect 62914 59726 62916 59778
rect 62860 59668 62916 59726
rect 62860 59612 63028 59668
rect 61628 59276 61796 59332
rect 61628 59106 61684 59118
rect 61628 59054 61630 59106
rect 61682 59054 61684 59106
rect 61628 58772 61684 59054
rect 61628 58210 61684 58716
rect 61628 58158 61630 58210
rect 61682 58158 61684 58210
rect 61628 57540 61684 58158
rect 61628 57474 61684 57484
rect 61516 56812 61684 56868
rect 61516 56644 61572 56654
rect 61404 56642 61572 56644
rect 61404 56590 61518 56642
rect 61570 56590 61572 56642
rect 61404 56588 61572 56590
rect 61516 56578 61572 56588
rect 60956 56252 61124 56308
rect 60844 56084 60900 56094
rect 60844 55990 60900 56028
rect 60620 55074 60676 55086
rect 60620 55022 60622 55074
rect 60674 55022 60676 55074
rect 60620 54852 60676 55022
rect 60620 54786 60676 54796
rect 60732 54402 60788 54414
rect 60732 54350 60734 54402
rect 60786 54350 60788 54402
rect 60732 53956 60788 54350
rect 60732 53890 60788 53900
rect 60508 53730 60564 53788
rect 60508 53678 60510 53730
rect 60562 53678 60564 53730
rect 60508 53666 60564 53678
rect 60060 53506 60228 53508
rect 60060 53454 60062 53506
rect 60114 53454 60228 53506
rect 60060 53452 60228 53454
rect 60060 53442 60116 53452
rect 60060 52834 60116 52846
rect 60060 52782 60062 52834
rect 60114 52782 60116 52834
rect 60060 52612 60116 52782
rect 60060 52546 60116 52556
rect 59948 51314 60004 51324
rect 59724 50594 59892 50596
rect 59724 50542 59726 50594
rect 59778 50542 59892 50594
rect 59724 50540 59892 50542
rect 59724 50530 59780 50540
rect 59276 50372 59444 50428
rect 58940 48850 58996 48860
rect 59052 49308 59220 49364
rect 58604 48738 58660 48748
rect 58156 48468 58212 48478
rect 58156 48354 58212 48412
rect 58156 48302 58158 48354
rect 58210 48302 58212 48354
rect 58156 48290 58212 48302
rect 58716 48466 58772 48478
rect 58716 48414 58718 48466
rect 58770 48414 58772 48466
rect 58380 48132 58436 48142
rect 58380 48038 58436 48076
rect 58604 48020 58660 48030
rect 58492 48018 58660 48020
rect 58492 47966 58606 48018
rect 58658 47966 58660 48018
rect 58492 47964 58660 47966
rect 58044 47852 58212 47908
rect 58156 46676 58212 47852
rect 58268 47684 58324 47694
rect 58492 47684 58548 47964
rect 58604 47954 58660 47964
rect 58268 47682 58548 47684
rect 58268 47630 58270 47682
rect 58322 47630 58548 47682
rect 58268 47628 58548 47630
rect 58716 47684 58772 48414
rect 58828 48356 58884 48366
rect 59052 48356 59108 49308
rect 59388 48468 59444 50372
rect 59500 50260 59556 50428
rect 59500 50194 59556 50204
rect 59388 48412 59780 48468
rect 58828 48354 59108 48356
rect 58828 48302 58830 48354
rect 58882 48302 59108 48354
rect 58828 48300 59108 48302
rect 58828 48290 58884 48300
rect 59164 48244 59220 48254
rect 59612 48244 59668 48254
rect 59164 48242 59668 48244
rect 59164 48190 59166 48242
rect 59218 48190 59614 48242
rect 59666 48190 59668 48242
rect 59164 48188 59668 48190
rect 59164 48178 59220 48188
rect 59612 48178 59668 48188
rect 58268 47618 58324 47628
rect 58716 47618 58772 47628
rect 59612 47684 59668 47694
rect 59612 47590 59668 47628
rect 59052 47460 59108 47470
rect 59052 47366 59108 47404
rect 58268 47348 58324 47358
rect 58268 46898 58324 47292
rect 58716 47346 58772 47358
rect 58716 47294 58718 47346
rect 58770 47294 58772 47346
rect 58716 47012 58772 47294
rect 58828 47348 58884 47358
rect 58828 47254 58884 47292
rect 58716 46946 58772 46956
rect 58268 46846 58270 46898
rect 58322 46846 58324 46898
rect 58268 46834 58324 46846
rect 57932 45826 57988 45836
rect 58044 46620 58156 46676
rect 56700 42868 56756 42878
rect 57148 42868 57204 45052
rect 57372 44434 57428 44446
rect 57372 44382 57374 44434
rect 57426 44382 57428 44434
rect 57260 42868 57316 42878
rect 56588 42866 56868 42868
rect 56588 42814 56702 42866
rect 56754 42814 56868 42866
rect 56588 42812 56868 42814
rect 57148 42866 57316 42868
rect 57148 42814 57262 42866
rect 57314 42814 57316 42866
rect 57148 42812 57316 42814
rect 56364 42774 56420 42812
rect 56700 42802 56756 42812
rect 55692 41970 55748 42588
rect 56812 42532 56868 42812
rect 57260 42802 57316 42812
rect 56812 42194 56868 42476
rect 56812 42142 56814 42194
rect 56866 42142 56868 42194
rect 56812 42130 56868 42142
rect 55692 41918 55694 41970
rect 55746 41918 55748 41970
rect 55692 41906 55748 41918
rect 56364 41972 56420 41982
rect 56364 41298 56420 41916
rect 57372 41858 57428 44382
rect 57820 43876 57876 45276
rect 58044 44100 58100 46620
rect 58156 46610 58212 46620
rect 59276 46674 59332 46686
rect 59276 46622 59278 46674
rect 59330 46622 59332 46674
rect 58604 46564 58660 46574
rect 58604 46470 58660 46508
rect 59276 46564 59332 46622
rect 58604 45892 58660 45902
rect 58604 45798 58660 45836
rect 58940 45892 58996 45902
rect 58940 45798 58996 45836
rect 58716 45666 58772 45678
rect 58716 45614 58718 45666
rect 58770 45614 58772 45666
rect 57820 43810 57876 43820
rect 57932 44044 58100 44100
rect 58268 45106 58324 45118
rect 58268 45054 58270 45106
rect 58322 45054 58324 45106
rect 57484 43652 57540 43662
rect 57484 43558 57540 43596
rect 57932 42868 57988 44044
rect 57932 42754 57988 42812
rect 57932 42702 57934 42754
rect 57986 42702 57988 42754
rect 57932 42690 57988 42702
rect 58044 43426 58100 43438
rect 58044 43374 58046 43426
rect 58098 43374 58100 43426
rect 58044 42756 58100 43374
rect 58268 42980 58324 45054
rect 58492 45108 58548 45118
rect 58492 45014 58548 45052
rect 58380 44994 58436 45006
rect 58380 44942 58382 44994
rect 58434 44942 58436 44994
rect 58380 44436 58436 44942
rect 58716 44996 58772 45614
rect 59276 45444 59332 46508
rect 59612 46114 59668 46126
rect 59612 46062 59614 46114
rect 59666 46062 59668 46114
rect 59612 45668 59668 46062
rect 59276 45378 59332 45388
rect 59388 45666 59668 45668
rect 59388 45614 59614 45666
rect 59666 45614 59668 45666
rect 59388 45612 59668 45614
rect 58828 45220 58884 45230
rect 58828 45126 58884 45164
rect 59388 45220 59444 45612
rect 59612 45602 59668 45612
rect 58380 44370 58436 44380
rect 58492 44884 58548 44894
rect 58492 43538 58548 44828
rect 58716 43708 58772 44940
rect 58492 43486 58494 43538
rect 58546 43486 58548 43538
rect 58268 42924 58436 42980
rect 58268 42756 58324 42766
rect 58044 42754 58324 42756
rect 58044 42702 58270 42754
rect 58322 42702 58324 42754
rect 58044 42700 58324 42702
rect 58268 42690 58324 42700
rect 57372 41806 57374 41858
rect 57426 41806 57428 41858
rect 56364 41246 56366 41298
rect 56418 41246 56420 41298
rect 56364 40740 56420 41246
rect 56364 40674 56420 40684
rect 57148 41410 57204 41422
rect 57148 41358 57150 41410
rect 57202 41358 57204 41410
rect 57148 41298 57204 41358
rect 57148 41246 57150 41298
rect 57202 41246 57204 41298
rect 55580 40226 55636 40236
rect 56476 40292 56532 40302
rect 56364 38162 56420 38174
rect 56364 38110 56366 38162
rect 56418 38110 56420 38162
rect 56028 37828 56084 37838
rect 56028 37490 56084 37772
rect 56364 37828 56420 38110
rect 56364 37762 56420 37772
rect 56028 37438 56030 37490
rect 56082 37438 56084 37490
rect 56028 37426 56084 37438
rect 56476 37268 56532 40236
rect 55468 37090 55524 37100
rect 56364 37156 56420 37166
rect 56476 37156 56532 37212
rect 56364 37154 56532 37156
rect 56364 37102 56366 37154
rect 56418 37102 56532 37154
rect 56364 37100 56532 37102
rect 54908 36978 54964 36988
rect 54796 20132 54964 20188
rect 54796 5012 54852 5022
rect 54796 4918 54852 4956
rect 54684 4174 54686 4226
rect 54738 4174 54740 4226
rect 54684 4162 54740 4174
rect 54684 3668 54740 3678
rect 54908 3668 54964 20132
rect 56364 9268 56420 37100
rect 57148 31108 57204 41246
rect 57372 41188 57428 41806
rect 57708 42642 57764 42654
rect 57708 42590 57710 42642
rect 57762 42590 57764 42642
rect 57708 41410 57764 42590
rect 58044 42530 58100 42542
rect 58044 42478 58046 42530
rect 58098 42478 58100 42530
rect 58044 42308 58100 42478
rect 58156 42532 58212 42542
rect 58380 42532 58436 42924
rect 58156 42438 58212 42476
rect 58268 42476 58436 42532
rect 58268 42308 58324 42476
rect 58044 42252 58324 42308
rect 58156 42084 58212 42094
rect 58156 41990 58212 42028
rect 57708 41358 57710 41410
rect 57762 41358 57764 41410
rect 57708 41346 57764 41358
rect 57932 41970 57988 41982
rect 57932 41918 57934 41970
rect 57986 41918 57988 41970
rect 57372 41122 57428 41132
rect 57596 40964 57652 40974
rect 57932 40964 57988 41918
rect 58268 41746 58324 41758
rect 58268 41694 58270 41746
rect 58322 41694 58324 41746
rect 58268 41300 58324 41694
rect 58268 41234 58324 41244
rect 58492 41188 58548 43486
rect 58492 41122 58548 41132
rect 58604 43652 58772 43708
rect 58940 45108 58996 45118
rect 57596 40962 57988 40964
rect 57596 40910 57598 40962
rect 57650 40910 57988 40962
rect 57596 40908 57988 40910
rect 58156 40962 58212 40974
rect 58156 40910 58158 40962
rect 58210 40910 58212 40962
rect 57596 39620 57652 40908
rect 57596 39554 57652 39564
rect 57708 40740 57764 40750
rect 57148 31042 57204 31052
rect 57708 34692 57764 40684
rect 58156 40628 58212 40910
rect 58156 40562 58212 40572
rect 58604 40292 58660 43652
rect 58940 43538 58996 45052
rect 58940 43486 58942 43538
rect 58994 43486 58996 43538
rect 58940 43474 58996 43486
rect 59276 45106 59332 45118
rect 59276 45054 59278 45106
rect 59330 45054 59332 45106
rect 59164 43316 59220 43326
rect 58716 42868 58772 42878
rect 58716 41298 58772 42812
rect 58716 41246 58718 41298
rect 58770 41246 58772 41298
rect 58716 41234 58772 41246
rect 58828 42866 58884 42878
rect 58828 42814 58830 42866
rect 58882 42814 58884 42866
rect 58828 40628 58884 42814
rect 59164 42754 59220 43260
rect 59164 42702 59166 42754
rect 59218 42702 59220 42754
rect 59164 42084 59220 42702
rect 59164 42018 59220 42028
rect 59276 41858 59332 45054
rect 59388 43652 59444 45164
rect 59500 45218 59556 45230
rect 59500 45166 59502 45218
rect 59554 45166 59556 45218
rect 59500 44884 59556 45166
rect 59612 45108 59668 45118
rect 59612 45014 59668 45052
rect 59500 44818 59556 44828
rect 59500 44436 59556 44446
rect 59500 44342 59556 44380
rect 59724 43764 59780 48412
rect 59836 47684 59892 50540
rect 59948 50596 60004 50606
rect 59948 50502 60004 50540
rect 59948 49026 60004 49038
rect 59948 48974 59950 49026
rect 60002 48974 60004 49026
rect 59948 48804 60004 48974
rect 60060 48916 60116 48926
rect 60060 48822 60116 48860
rect 59948 48738 60004 48748
rect 59836 47618 59892 47628
rect 59948 47570 60004 47582
rect 59948 47518 59950 47570
rect 60002 47518 60004 47570
rect 59836 47234 59892 47246
rect 59836 47182 59838 47234
rect 59890 47182 59892 47234
rect 59836 46114 59892 47182
rect 59948 46786 60004 47518
rect 59948 46734 59950 46786
rect 60002 46734 60004 46786
rect 59948 46722 60004 46734
rect 59836 46062 59838 46114
rect 59890 46062 59892 46114
rect 59836 46050 59892 46062
rect 60172 45892 60228 53452
rect 60956 53284 61012 56252
rect 61292 56082 61348 56094
rect 61292 56030 61294 56082
rect 61346 56030 61348 56082
rect 61292 55412 61348 56030
rect 61292 55410 61460 55412
rect 61292 55358 61294 55410
rect 61346 55358 61460 55410
rect 61292 55356 61460 55358
rect 61292 55346 61348 55356
rect 60620 53228 61012 53284
rect 61292 53954 61348 53966
rect 61292 53902 61294 53954
rect 61346 53902 61348 53954
rect 61292 53506 61348 53902
rect 61404 53732 61460 55356
rect 61404 53666 61460 53676
rect 61292 53454 61294 53506
rect 61346 53454 61348 53506
rect 60508 53060 60564 53070
rect 60508 52966 60564 53004
rect 60620 52612 60676 53228
rect 61292 53172 61348 53454
rect 61628 53284 61684 56812
rect 61740 56420 61796 59276
rect 62076 59220 62132 59230
rect 62076 59126 62132 59164
rect 62188 58772 62244 58782
rect 62188 58658 62244 58716
rect 62188 58606 62190 58658
rect 62242 58606 62244 58658
rect 62188 58594 62244 58606
rect 62524 58660 62580 58670
rect 62636 58660 62692 59500
rect 62860 59444 62916 59454
rect 62860 59350 62916 59388
rect 62748 59220 62804 59230
rect 62748 59126 62804 59164
rect 62972 59108 63028 59612
rect 63084 59218 63140 60174
rect 63084 59166 63086 59218
rect 63138 59166 63140 59218
rect 63084 59154 63140 59166
rect 62524 58658 62692 58660
rect 62524 58606 62526 58658
rect 62578 58606 62692 58658
rect 62524 58604 62692 58606
rect 62860 58884 62916 58894
rect 62524 58594 62580 58604
rect 62412 58210 62468 58222
rect 62412 58158 62414 58210
rect 62466 58158 62468 58210
rect 62412 57876 62468 58158
rect 62412 57810 62468 57820
rect 62860 57874 62916 58828
rect 62860 57822 62862 57874
rect 62914 57822 62916 57874
rect 62860 57810 62916 57822
rect 61964 57764 62020 57774
rect 61852 57540 61908 57550
rect 61852 57446 61908 57484
rect 61964 56978 62020 57708
rect 61964 56926 61966 56978
rect 62018 56926 62020 56978
rect 61964 56914 62020 56926
rect 62300 57650 62356 57662
rect 62972 57652 63028 59052
rect 63084 58548 63140 58558
rect 63196 58548 63252 61628
rect 63308 59890 63364 59902
rect 63308 59838 63310 59890
rect 63362 59838 63364 59890
rect 63308 59330 63364 59838
rect 63308 59278 63310 59330
rect 63362 59278 63364 59330
rect 63308 59266 63364 59278
rect 63084 58546 63252 58548
rect 63084 58494 63086 58546
rect 63138 58494 63252 58546
rect 63084 58492 63252 58494
rect 63084 58482 63140 58492
rect 62300 57598 62302 57650
rect 62354 57598 62356 57650
rect 62300 56980 62356 57598
rect 62748 57596 63028 57652
rect 62300 56532 62356 56924
rect 62636 56980 62692 56990
rect 62524 56756 62580 56766
rect 62636 56756 62692 56924
rect 62580 56700 62692 56756
rect 62524 56690 62580 56700
rect 62300 56466 62356 56476
rect 61740 56364 62020 56420
rect 61740 55970 61796 55982
rect 61740 55918 61742 55970
rect 61794 55918 61796 55970
rect 61740 55300 61796 55918
rect 61740 55234 61796 55244
rect 61852 55298 61908 55310
rect 61852 55246 61854 55298
rect 61906 55246 61908 55298
rect 61740 54292 61796 54302
rect 61740 53730 61796 54236
rect 61852 53954 61908 55246
rect 61852 53902 61854 53954
rect 61906 53902 61908 53954
rect 61852 53890 61908 53902
rect 61740 53678 61742 53730
rect 61794 53678 61796 53730
rect 61740 53666 61796 53678
rect 61852 53284 61908 53294
rect 61628 53228 61796 53284
rect 60844 53116 61348 53172
rect 60508 52556 60676 52612
rect 60732 52722 60788 52734
rect 60732 52670 60734 52722
rect 60786 52670 60788 52722
rect 60284 52388 60340 52398
rect 60284 52294 60340 52332
rect 60508 52164 60564 52556
rect 60620 52388 60676 52398
rect 60732 52388 60788 52670
rect 60620 52386 60788 52388
rect 60620 52334 60622 52386
rect 60674 52334 60788 52386
rect 60620 52332 60788 52334
rect 60620 52322 60676 52332
rect 60396 52108 60564 52164
rect 60396 51828 60452 52108
rect 60508 51940 60564 51950
rect 60508 51938 60788 51940
rect 60508 51886 60510 51938
rect 60562 51886 60788 51938
rect 60508 51884 60788 51886
rect 60508 51874 60564 51884
rect 60284 51380 60340 51390
rect 60284 51286 60340 51324
rect 60396 50708 60452 51772
rect 60620 51380 60676 51390
rect 60508 50708 60564 50718
rect 60396 50706 60564 50708
rect 60396 50654 60510 50706
rect 60562 50654 60564 50706
rect 60396 50652 60564 50654
rect 60508 50642 60564 50652
rect 60620 49922 60676 51324
rect 60620 49870 60622 49922
rect 60674 49870 60676 49922
rect 60620 49858 60676 49870
rect 60620 49364 60676 49374
rect 60060 45836 60228 45892
rect 60284 49140 60340 49150
rect 60060 45220 60116 45836
rect 60172 45668 60228 45678
rect 60284 45668 60340 49084
rect 60620 48804 60676 49308
rect 60732 49028 60788 51884
rect 60732 48962 60788 48972
rect 60508 48242 60564 48254
rect 60508 48190 60510 48242
rect 60562 48190 60564 48242
rect 60396 48132 60452 48142
rect 60396 48038 60452 48076
rect 60172 45666 60340 45668
rect 60172 45614 60174 45666
rect 60226 45614 60340 45666
rect 60172 45612 60340 45614
rect 60396 47684 60452 47694
rect 60396 47570 60452 47628
rect 60396 47518 60398 47570
rect 60450 47518 60452 47570
rect 60172 45602 60228 45612
rect 60284 45444 60340 45454
rect 60060 45164 60228 45220
rect 60060 44994 60116 45006
rect 60060 44942 60062 44994
rect 60114 44942 60116 44994
rect 60060 44884 60116 44942
rect 60060 44100 60116 44828
rect 60060 44034 60116 44044
rect 59948 43764 60004 43774
rect 59724 43762 60004 43764
rect 59724 43710 59950 43762
rect 60002 43710 60004 43762
rect 59724 43708 60004 43710
rect 59948 43698 60004 43708
rect 59388 43586 59444 43596
rect 59612 43540 59668 43550
rect 60172 43540 60228 45164
rect 60284 44322 60340 45388
rect 60284 44270 60286 44322
rect 60338 44270 60340 44322
rect 60284 44258 60340 44270
rect 59612 42754 59668 43484
rect 59612 42702 59614 42754
rect 59666 42702 59668 42754
rect 59388 42644 59444 42654
rect 59388 42530 59444 42588
rect 59388 42478 59390 42530
rect 59442 42478 59444 42530
rect 59388 42466 59444 42478
rect 59500 42642 59556 42654
rect 59500 42590 59502 42642
rect 59554 42590 59556 42642
rect 59388 42084 59444 42094
rect 59388 41970 59444 42028
rect 59388 41918 59390 41970
rect 59442 41918 59444 41970
rect 59388 41906 59444 41918
rect 59276 41806 59278 41858
rect 59330 41806 59332 41858
rect 59276 41794 59332 41806
rect 59500 41746 59556 42590
rect 59612 42532 59668 42702
rect 59836 43484 60228 43540
rect 60284 43764 60340 43774
rect 60284 43538 60340 43708
rect 60284 43486 60286 43538
rect 60338 43486 60340 43538
rect 59836 42532 59892 43484
rect 60284 43474 60340 43486
rect 59948 43316 60004 43326
rect 59948 43222 60004 43260
rect 60060 43314 60116 43326
rect 60060 43262 60062 43314
rect 60114 43262 60116 43314
rect 60060 43092 60116 43262
rect 60060 43026 60116 43036
rect 59948 42868 60004 42878
rect 59948 42754 60004 42812
rect 59948 42702 59950 42754
rect 60002 42702 60004 42754
rect 59948 42690 60004 42702
rect 59836 42476 60004 42532
rect 59612 42466 59668 42476
rect 59500 41694 59502 41746
rect 59554 41694 59556 41746
rect 59500 41682 59556 41694
rect 59836 41972 59892 41982
rect 59500 41300 59556 41310
rect 59500 41206 59556 41244
rect 59052 41188 59108 41198
rect 59052 41094 59108 41132
rect 58828 40562 58884 40572
rect 58604 40226 58660 40236
rect 58268 34802 58324 34814
rect 58268 34750 58270 34802
rect 58322 34750 58324 34802
rect 58268 34692 58324 34750
rect 57708 34690 58324 34692
rect 57708 34638 57710 34690
rect 57762 34638 58324 34690
rect 57708 34636 58324 34638
rect 58604 34692 58660 34702
rect 56364 9202 56420 9212
rect 57708 8428 57764 34636
rect 58604 34598 58660 34636
rect 58828 32004 58884 32014
rect 58828 26402 58884 31948
rect 58828 26350 58830 26402
rect 58882 26350 58884 26402
rect 58828 26338 58884 26350
rect 59836 22260 59892 41916
rect 59836 22194 59892 22204
rect 57372 8372 57764 8428
rect 55244 5012 55300 5022
rect 55244 4918 55300 4956
rect 57372 4562 57428 8372
rect 59948 6020 60004 42476
rect 60060 42530 60116 42542
rect 60060 42478 60062 42530
rect 60114 42478 60116 42530
rect 60060 41746 60116 42478
rect 60060 41694 60062 41746
rect 60114 41694 60116 41746
rect 60060 41682 60116 41694
rect 60172 42084 60228 42094
rect 60396 42084 60452 47518
rect 60508 45444 60564 48190
rect 60620 46002 60676 48748
rect 60844 46788 60900 53116
rect 61404 52948 61460 52958
rect 61404 52854 61460 52892
rect 60956 52834 61012 52846
rect 60956 52782 60958 52834
rect 61010 52782 61012 52834
rect 60956 52388 61012 52782
rect 60956 52322 61012 52332
rect 61404 52722 61460 52734
rect 61404 52670 61406 52722
rect 61458 52670 61460 52722
rect 61404 52162 61460 52670
rect 61404 52110 61406 52162
rect 61458 52110 61460 52162
rect 61404 52098 61460 52110
rect 61516 52388 61572 52398
rect 61068 51266 61124 51278
rect 61068 51214 61070 51266
rect 61122 51214 61124 51266
rect 61068 50428 61124 51214
rect 61516 50818 61572 52332
rect 61516 50766 61518 50818
rect 61570 50766 61572 50818
rect 61068 50372 61460 50428
rect 61292 49700 61348 49710
rect 60844 46722 60900 46732
rect 61068 49476 61124 49486
rect 60620 45950 60622 46002
rect 60674 45950 60676 46002
rect 60620 45938 60676 45950
rect 60844 46228 60900 46238
rect 60508 45388 60676 45444
rect 60508 44994 60564 45006
rect 60508 44942 60510 44994
rect 60562 44942 60564 44994
rect 60508 43540 60564 44942
rect 60620 44882 60676 45388
rect 60620 44830 60622 44882
rect 60674 44830 60676 44882
rect 60620 44818 60676 44830
rect 60508 43474 60564 43484
rect 60508 43314 60564 43326
rect 60508 43262 60510 43314
rect 60562 43262 60564 43314
rect 60508 42980 60564 43262
rect 60844 43316 60900 46172
rect 60956 44994 61012 45006
rect 60956 44942 60958 44994
rect 61010 44942 61012 44994
rect 60956 44882 61012 44942
rect 60956 44830 60958 44882
rect 61010 44830 61012 44882
rect 60956 43540 61012 44830
rect 61068 44660 61124 49420
rect 61180 48916 61236 48926
rect 61292 48916 61348 49644
rect 61404 49140 61460 50372
rect 61516 49364 61572 50766
rect 61628 50708 61684 50718
rect 61628 50484 61684 50652
rect 61628 50418 61684 50428
rect 61516 49298 61572 49308
rect 61516 49140 61572 49150
rect 61404 49138 61572 49140
rect 61404 49086 61518 49138
rect 61570 49086 61572 49138
rect 61404 49084 61572 49086
rect 61516 49074 61572 49084
rect 61740 49140 61796 53228
rect 61852 53170 61908 53228
rect 61852 53118 61854 53170
rect 61906 53118 61908 53170
rect 61852 52500 61908 53118
rect 61852 52434 61908 52444
rect 61628 49028 61684 49038
rect 61628 48934 61684 48972
rect 61404 48916 61460 48926
rect 61292 48914 61460 48916
rect 61292 48862 61406 48914
rect 61458 48862 61460 48914
rect 61292 48860 61460 48862
rect 61180 47460 61236 48860
rect 61404 48850 61460 48860
rect 61740 48692 61796 49084
rect 61628 48636 61796 48692
rect 61292 48242 61348 48254
rect 61292 48190 61294 48242
rect 61346 48190 61348 48242
rect 61292 47908 61348 48190
rect 61516 48244 61572 48254
rect 61516 48150 61572 48188
rect 61404 48132 61460 48142
rect 61404 48038 61460 48076
rect 61292 47842 61348 47852
rect 61292 47460 61348 47470
rect 61180 47458 61348 47460
rect 61180 47406 61294 47458
rect 61346 47406 61348 47458
rect 61180 47404 61348 47406
rect 61292 47394 61348 47404
rect 61628 47458 61684 48636
rect 61740 48356 61796 48366
rect 61740 48262 61796 48300
rect 61628 47406 61630 47458
rect 61682 47406 61684 47458
rect 61628 47394 61684 47406
rect 61852 48132 61908 48142
rect 61852 47908 61908 48076
rect 61516 47234 61572 47246
rect 61516 47182 61518 47234
rect 61570 47182 61572 47234
rect 61404 45890 61460 45902
rect 61404 45838 61406 45890
rect 61458 45838 61460 45890
rect 61404 45332 61460 45838
rect 61516 45332 61572 47182
rect 61628 45332 61684 45342
rect 61516 45330 61684 45332
rect 61516 45278 61630 45330
rect 61682 45278 61684 45330
rect 61516 45276 61684 45278
rect 61404 45266 61460 45276
rect 61068 44594 61124 44604
rect 61292 45108 61348 45118
rect 61292 44324 61348 45052
rect 61628 44436 61684 45276
rect 61852 45332 61908 47852
rect 61964 46564 62020 56364
rect 62412 56308 62468 56318
rect 62188 56252 62412 56308
rect 62076 55412 62132 55422
rect 62076 55318 62132 55356
rect 62188 53844 62244 56252
rect 62412 56214 62468 56252
rect 62300 55300 62356 55338
rect 62300 55234 62356 55244
rect 62524 55298 62580 55310
rect 62524 55246 62526 55298
rect 62578 55246 62580 55298
rect 62300 55076 62356 55086
rect 62300 54982 62356 55020
rect 62188 53788 62356 53844
rect 62188 53620 62244 53630
rect 62188 53526 62244 53564
rect 62076 53172 62132 53182
rect 62076 52836 62132 53116
rect 62300 53060 62356 53788
rect 62076 52770 62132 52780
rect 62188 53004 62356 53060
rect 62524 53508 62580 55246
rect 62748 54404 62804 57596
rect 63308 57538 63364 57550
rect 63308 57486 63310 57538
rect 63362 57486 63364 57538
rect 63308 56980 63364 57486
rect 63308 56914 63364 56924
rect 62860 55972 62916 55982
rect 62860 55878 62916 55916
rect 62860 55300 62916 55310
rect 62860 54964 62916 55244
rect 62972 55188 63028 55198
rect 62972 55094 63028 55132
rect 62860 54898 62916 54908
rect 63196 54628 63252 54638
rect 62748 54338 62804 54348
rect 62972 54404 63028 54414
rect 62972 54310 63028 54348
rect 62188 51940 62244 53004
rect 62300 52834 62356 52846
rect 62300 52782 62302 52834
rect 62354 52782 62356 52834
rect 62300 52052 62356 52782
rect 62524 52500 62580 53452
rect 62524 52434 62580 52444
rect 62636 53732 62692 53742
rect 62300 51986 62356 51996
rect 62412 52388 62468 52398
rect 62188 51874 62244 51884
rect 62076 50820 62132 50830
rect 62076 49026 62132 50764
rect 62076 48974 62078 49026
rect 62130 48974 62132 49026
rect 62076 48962 62132 48974
rect 62188 50596 62244 50606
rect 62188 47682 62244 50540
rect 62412 50428 62468 52332
rect 62636 51380 62692 53676
rect 63084 52612 63140 52622
rect 63084 52274 63140 52556
rect 63084 52222 63086 52274
rect 63138 52222 63140 52274
rect 63084 52210 63140 52222
rect 62636 51314 62692 51324
rect 63084 51940 63140 51950
rect 62412 50372 62580 50428
rect 62524 49140 62580 50372
rect 62860 49700 62916 49710
rect 62524 49084 62692 49140
rect 62188 47630 62190 47682
rect 62242 47630 62244 47682
rect 62188 47618 62244 47630
rect 62412 48916 62468 48926
rect 62412 47572 62468 48860
rect 62524 48244 62580 48254
rect 62524 47796 62580 48188
rect 62524 47730 62580 47740
rect 62636 47684 62692 49084
rect 62860 49026 62916 49644
rect 62972 49140 63028 49150
rect 62972 49046 63028 49084
rect 62860 48974 62862 49026
rect 62914 48974 62916 49026
rect 62748 48802 62804 48814
rect 62748 48750 62750 48802
rect 62802 48750 62804 48802
rect 62748 48020 62804 48750
rect 62860 48244 62916 48974
rect 63084 48916 63140 51884
rect 63196 50708 63252 54572
rect 63308 53732 63364 53742
rect 63308 53638 63364 53676
rect 63308 52836 63364 52846
rect 63308 52742 63364 52780
rect 63420 52388 63476 62132
rect 63532 60786 63588 60798
rect 63532 60734 63534 60786
rect 63586 60734 63588 60786
rect 63532 60116 63588 60734
rect 63756 60674 63812 62300
rect 63756 60622 63758 60674
rect 63810 60622 63812 60674
rect 63756 60610 63812 60622
rect 63868 62354 63924 62366
rect 63868 62302 63870 62354
rect 63922 62302 63924 62354
rect 63532 60022 63588 60060
rect 63644 60564 63700 60574
rect 63644 59442 63700 60508
rect 63868 60116 63924 62302
rect 64092 62354 64148 62524
rect 64652 62514 64708 62524
rect 64092 62302 64094 62354
rect 64146 62302 64148 62354
rect 64092 62290 64148 62302
rect 64876 62188 64932 63980
rect 64428 62132 64932 62188
rect 64428 60674 64484 62132
rect 64988 60788 65044 65548
rect 65212 62188 65268 114268
rect 65916 113708 66180 113718
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 65916 113642 66180 113652
rect 67788 113428 67844 113438
rect 65916 112140 66180 112150
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 65916 112074 66180 112084
rect 65916 110572 66180 110582
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 65916 110506 66180 110516
rect 65916 109004 66180 109014
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 65916 108938 66180 108948
rect 65916 107436 66180 107446
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 65916 107370 66180 107380
rect 65916 105868 66180 105878
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 65916 105802 66180 105812
rect 65916 104300 66180 104310
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 65916 104234 66180 104244
rect 65916 102732 66180 102742
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 65916 102666 66180 102676
rect 65916 101164 66180 101174
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 65916 101098 66180 101108
rect 65916 99596 66180 99606
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 65916 99530 66180 99540
rect 65916 98028 66180 98038
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 65916 97962 66180 97972
rect 65916 96460 66180 96470
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 65916 96394 66180 96404
rect 65916 94892 66180 94902
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 65916 94826 66180 94836
rect 65916 93324 66180 93334
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 65916 93258 66180 93268
rect 65916 91756 66180 91766
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 65916 91690 66180 91700
rect 65916 90188 66180 90198
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 65916 90122 66180 90132
rect 65916 88620 66180 88630
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 65916 88554 66180 88564
rect 65916 87052 66180 87062
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 65916 86986 66180 86996
rect 65916 85484 66180 85494
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 65916 85418 66180 85428
rect 65916 83916 66180 83926
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 65916 83850 66180 83860
rect 65916 82348 66180 82358
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 65916 82282 66180 82292
rect 65916 80780 66180 80790
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 65916 80714 66180 80724
rect 65916 79212 66180 79222
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 65916 79146 66180 79156
rect 65916 77644 66180 77654
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 65916 77578 66180 77588
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 67340 68068 67396 68078
rect 65324 67060 65380 67070
rect 65324 66966 65380 67004
rect 65660 67060 65716 67070
rect 65324 66052 65380 66062
rect 65324 64706 65380 65996
rect 65660 65604 65716 67004
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65884 66386 65940 66398
rect 65884 66334 65886 66386
rect 65938 66334 65940 66386
rect 65884 66052 65940 66334
rect 67116 66164 67172 66174
rect 65884 65986 65940 65996
rect 66332 66052 66388 66062
rect 66332 65958 66388 65996
rect 66780 66050 66836 66062
rect 66780 65998 66782 66050
rect 66834 65998 66836 66050
rect 65660 65490 65716 65548
rect 65660 65438 65662 65490
rect 65714 65438 65716 65490
rect 65660 65426 65716 65438
rect 66780 65604 66836 65998
rect 66444 65380 66500 65390
rect 66332 65378 66500 65380
rect 66332 65326 66446 65378
rect 66498 65326 66500 65378
rect 66332 65324 66500 65326
rect 65324 64654 65326 64706
rect 65378 64654 65380 64706
rect 65324 64642 65380 64654
rect 65772 65268 65828 65278
rect 65772 64708 65828 65212
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 65996 64708 66052 64718
rect 65772 64652 65996 64708
rect 65996 64576 66052 64652
rect 65436 64484 65492 64494
rect 65436 64390 65492 64428
rect 66332 64482 66388 65324
rect 66444 65314 66500 65324
rect 66332 64430 66334 64482
rect 66386 64430 66388 64482
rect 66332 64418 66388 64430
rect 66444 64594 66500 64606
rect 66444 64542 66446 64594
rect 66498 64542 66500 64594
rect 66444 64484 66500 64542
rect 65548 64372 65604 64382
rect 65548 64146 65604 64316
rect 65548 64094 65550 64146
rect 65602 64094 65604 64146
rect 65548 64082 65604 64094
rect 65660 64036 65716 64046
rect 65660 63942 65716 63980
rect 65324 63924 65380 63934
rect 65324 63830 65380 63868
rect 65548 63812 65604 63822
rect 65548 63588 65604 63756
rect 66220 63812 66276 63822
rect 66276 63756 66388 63812
rect 66220 63718 66276 63756
rect 66332 63588 66388 63756
rect 65436 63140 65492 63150
rect 65548 63140 65604 63532
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66332 63522 66388 63532
rect 65916 63466 66180 63476
rect 65436 63138 65604 63140
rect 65436 63086 65438 63138
rect 65490 63086 65604 63138
rect 65436 63084 65604 63086
rect 65436 63074 65492 63084
rect 65436 62916 65492 62926
rect 65436 62356 65492 62860
rect 64988 60722 65044 60732
rect 65100 62132 65268 62188
rect 65324 62354 65492 62356
rect 65324 62302 65438 62354
rect 65490 62302 65492 62354
rect 65324 62300 65492 62302
rect 64428 60622 64430 60674
rect 64482 60622 64484 60674
rect 63868 60050 63924 60060
rect 64092 60452 64148 60462
rect 63644 59390 63646 59442
rect 63698 59390 63700 59442
rect 63644 59378 63700 59390
rect 63532 59108 63588 59118
rect 63532 59014 63588 59052
rect 63980 59108 64036 59118
rect 63980 59014 64036 59052
rect 63980 58660 64036 58670
rect 64092 58660 64148 60396
rect 64428 60116 64484 60622
rect 64876 60676 64932 60686
rect 64876 60564 64932 60620
rect 64876 60508 65044 60564
rect 64316 59444 64372 59454
rect 64428 59444 64484 60060
rect 64316 59442 64484 59444
rect 64316 59390 64318 59442
rect 64370 59390 64484 59442
rect 64316 59388 64484 59390
rect 64316 59378 64372 59388
rect 64764 58884 64820 58894
rect 64204 58660 64260 58670
rect 63980 58658 64260 58660
rect 63980 58606 63982 58658
rect 64034 58606 64206 58658
rect 64258 58606 64260 58658
rect 63980 58604 64260 58606
rect 63980 58594 64036 58604
rect 64204 58594 64260 58604
rect 63644 58546 63700 58558
rect 63644 58494 63646 58546
rect 63698 58494 63700 58546
rect 63644 57650 63700 58494
rect 63756 58324 63812 58334
rect 63756 58230 63812 58268
rect 64540 58210 64596 58222
rect 64540 58158 64542 58210
rect 64594 58158 64596 58210
rect 64540 57876 64596 58158
rect 63980 57820 64372 57876
rect 63980 57762 64036 57820
rect 63980 57710 63982 57762
rect 64034 57710 64036 57762
rect 63980 57698 64036 57710
rect 63644 57598 63646 57650
rect 63698 57598 63700 57650
rect 63644 57586 63700 57598
rect 64092 57650 64148 57662
rect 64092 57598 64094 57650
rect 64146 57598 64148 57650
rect 63532 57538 63588 57550
rect 63532 57486 63534 57538
rect 63586 57486 63588 57538
rect 63532 57092 63588 57486
rect 63532 57026 63588 57036
rect 63980 56980 64036 56990
rect 63980 56866 64036 56924
rect 63980 56814 63982 56866
rect 64034 56814 64036 56866
rect 63532 56532 63588 56542
rect 63532 56194 63588 56476
rect 63532 56142 63534 56194
rect 63586 56142 63588 56194
rect 63532 56130 63588 56142
rect 63756 56196 63812 56234
rect 63756 56130 63812 56140
rect 63644 55970 63700 55982
rect 63644 55918 63646 55970
rect 63698 55918 63700 55970
rect 63644 55412 63700 55918
rect 63644 55346 63700 55356
rect 63756 55972 63812 55982
rect 63532 55074 63588 55086
rect 63532 55022 63534 55074
rect 63586 55022 63588 55074
rect 63532 53508 63588 55022
rect 63644 55076 63700 55086
rect 63644 54626 63700 55020
rect 63644 54574 63646 54626
rect 63698 54574 63700 54626
rect 63644 54562 63700 54574
rect 63756 54404 63812 55916
rect 63980 55524 64036 56814
rect 64092 56308 64148 57598
rect 64316 57092 64372 57820
rect 64540 57810 64596 57820
rect 64428 57650 64484 57662
rect 64428 57598 64430 57650
rect 64482 57598 64484 57650
rect 64428 57428 64484 57598
rect 64652 57650 64708 57662
rect 64652 57598 64654 57650
rect 64706 57598 64708 57650
rect 64652 57540 64708 57598
rect 64652 57474 64708 57484
rect 64428 57372 64596 57428
rect 64316 57036 64484 57092
rect 64428 56978 64484 57036
rect 64428 56926 64430 56978
rect 64482 56926 64484 56978
rect 64428 56914 64484 56926
rect 64316 56868 64372 56878
rect 64316 56774 64372 56812
rect 64092 56242 64148 56252
rect 64316 56532 64372 56542
rect 64316 56306 64372 56476
rect 64316 56254 64318 56306
rect 64370 56254 64372 56306
rect 63980 55458 64036 55468
rect 64204 56196 64260 56206
rect 64204 55410 64260 56140
rect 64204 55358 64206 55410
rect 64258 55358 64260 55410
rect 64204 55346 64260 55358
rect 63532 53442 63588 53452
rect 63644 54348 63812 54404
rect 63868 54740 63924 54750
rect 63868 54626 63924 54684
rect 63868 54574 63870 54626
rect 63922 54574 63924 54626
rect 63420 52322 63476 52332
rect 63196 50034 63252 50652
rect 63196 49982 63198 50034
rect 63250 49982 63252 50034
rect 63196 49970 63252 49982
rect 63308 51266 63364 51278
rect 63308 51214 63310 51266
rect 63362 51214 63364 51266
rect 63084 48850 63140 48860
rect 63196 49026 63252 49038
rect 63196 48974 63198 49026
rect 63250 48974 63252 49026
rect 62860 48178 62916 48188
rect 63084 48692 63140 48702
rect 63084 48356 63140 48636
rect 63084 48242 63140 48300
rect 63084 48190 63086 48242
rect 63138 48190 63140 48242
rect 63084 48178 63140 48190
rect 63084 48020 63140 48030
rect 62748 47964 63084 48020
rect 62972 47684 63028 47694
rect 62636 47628 62804 47684
rect 62412 47516 62692 47572
rect 62300 47458 62356 47470
rect 62300 47406 62302 47458
rect 62354 47406 62356 47458
rect 62300 46900 62356 47406
rect 62300 46834 62356 46844
rect 62636 46786 62692 47516
rect 62636 46734 62638 46786
rect 62690 46734 62692 46786
rect 62636 46722 62692 46734
rect 62076 46564 62132 46574
rect 61964 46562 62132 46564
rect 61964 46510 62078 46562
rect 62130 46510 62132 46562
rect 61964 46508 62132 46510
rect 61964 45332 62020 45342
rect 61852 45330 62020 45332
rect 61852 45278 61966 45330
rect 62018 45278 62020 45330
rect 61852 45276 62020 45278
rect 61628 44370 61684 44380
rect 61740 44996 61796 45006
rect 61292 44322 61572 44324
rect 61292 44270 61294 44322
rect 61346 44270 61572 44322
rect 61292 44268 61572 44270
rect 61292 44258 61348 44268
rect 61516 44212 61572 44268
rect 61516 43764 61572 44156
rect 61628 44100 61684 44110
rect 61628 44006 61684 44044
rect 61628 43764 61684 43774
rect 61516 43762 61684 43764
rect 61516 43710 61630 43762
rect 61682 43710 61684 43762
rect 61516 43708 61684 43710
rect 61628 43698 61684 43708
rect 61740 43652 61796 44940
rect 61852 44324 61908 45276
rect 61964 45266 62020 45276
rect 62076 44882 62132 46508
rect 62748 45220 62804 47628
rect 62972 47590 63028 47628
rect 63084 47570 63140 47964
rect 63196 48018 63252 48974
rect 63308 48468 63364 51214
rect 63644 50428 63700 54348
rect 63868 53732 63924 54574
rect 64316 54516 64372 56254
rect 64540 55972 64596 57372
rect 64540 55906 64596 55916
rect 64652 55524 64708 55534
rect 64652 55410 64708 55468
rect 64652 55358 64654 55410
rect 64706 55358 64708 55410
rect 64652 55346 64708 55358
rect 64428 54740 64484 54778
rect 64764 54740 64820 58828
rect 64876 58324 64932 58334
rect 64876 58230 64932 58268
rect 64988 56980 65044 60508
rect 64988 56914 65044 56924
rect 64484 54684 64820 54740
rect 64876 55636 64932 55646
rect 64428 54674 64484 54684
rect 64204 54460 64372 54516
rect 63980 54290 64036 54302
rect 63980 54238 63982 54290
rect 64034 54238 64036 54290
rect 63980 53842 64036 54238
rect 63980 53790 63982 53842
rect 64034 53790 64036 53842
rect 63980 53778 64036 53790
rect 63756 53676 63924 53732
rect 63756 52836 63812 53676
rect 64204 53172 64260 54460
rect 64204 53106 64260 53116
rect 63868 52948 63924 52958
rect 63868 52946 64036 52948
rect 63868 52894 63870 52946
rect 63922 52894 64036 52946
rect 63868 52892 64036 52894
rect 63868 52882 63924 52892
rect 63756 52770 63812 52780
rect 63980 52164 64036 52892
rect 64540 52834 64596 52846
rect 64540 52782 64542 52834
rect 64594 52782 64596 52834
rect 64428 52276 64484 52286
rect 64428 52182 64484 52220
rect 64540 52164 64596 52782
rect 63980 52162 64148 52164
rect 63980 52110 63982 52162
rect 64034 52110 64148 52162
rect 63980 52108 64148 52110
rect 63980 52098 64036 52108
rect 63868 51380 63924 51390
rect 63756 50708 63812 50718
rect 63756 50594 63812 50652
rect 63756 50542 63758 50594
rect 63810 50542 63812 50594
rect 63756 50530 63812 50542
rect 63420 50370 63476 50382
rect 63420 50318 63422 50370
rect 63474 50318 63476 50370
rect 63420 49924 63476 50318
rect 63420 49028 63476 49868
rect 63420 48962 63476 48972
rect 63532 50372 63700 50428
rect 63308 48412 63476 48468
rect 63308 48244 63364 48254
rect 63308 48150 63364 48188
rect 63420 48132 63476 48412
rect 63420 48066 63476 48076
rect 63196 47966 63198 48018
rect 63250 47966 63252 48018
rect 63196 47954 63252 47966
rect 63084 47518 63086 47570
rect 63138 47518 63140 47570
rect 63084 47506 63140 47518
rect 63308 47458 63364 47470
rect 63308 47406 63310 47458
rect 63362 47406 63364 47458
rect 63196 46788 63252 46798
rect 63196 46694 63252 46732
rect 62860 46674 62916 46686
rect 62860 46622 62862 46674
rect 62914 46622 62916 46674
rect 62860 46004 62916 46622
rect 62972 46676 63028 46686
rect 62972 46582 63028 46620
rect 63084 46674 63140 46686
rect 63084 46622 63086 46674
rect 63138 46622 63140 46674
rect 63084 46564 63140 46622
rect 63084 46498 63140 46508
rect 62860 45948 63028 46004
rect 62076 44830 62078 44882
rect 62130 44830 62132 44882
rect 62076 44818 62132 44830
rect 62636 45164 62804 45220
rect 62860 45780 62916 45790
rect 62860 45444 62916 45724
rect 61964 44548 62020 44558
rect 61964 44454 62020 44492
rect 62188 44324 62244 44334
rect 61852 44268 62020 44324
rect 61180 43540 61236 43550
rect 61740 43540 61796 43596
rect 60956 43484 61180 43540
rect 60844 43260 61124 43316
rect 60508 42914 60564 42924
rect 60620 43092 60676 43102
rect 60620 42866 60676 43036
rect 60620 42814 60622 42866
rect 60674 42814 60676 42866
rect 60620 42802 60676 42814
rect 60172 40964 60228 42028
rect 60284 42028 60452 42084
rect 60284 41300 60340 42028
rect 60956 41970 61012 41982
rect 60956 41918 60958 41970
rect 61010 41918 61012 41970
rect 60284 41234 60340 41244
rect 60396 41858 60452 41870
rect 60396 41806 60398 41858
rect 60450 41806 60452 41858
rect 60396 41746 60452 41806
rect 60396 41694 60398 41746
rect 60450 41694 60452 41746
rect 60172 40962 60340 40964
rect 60172 40910 60174 40962
rect 60226 40910 60340 40962
rect 60172 40908 60340 40910
rect 60172 40898 60228 40908
rect 60284 33012 60340 40908
rect 60172 32956 60340 33012
rect 59948 5954 60004 5964
rect 60060 32788 60116 32798
rect 57372 4510 57374 4562
rect 57426 4510 57428 4562
rect 56588 4340 56644 4350
rect 56588 4246 56644 4284
rect 57372 4340 57428 4510
rect 59836 5122 59892 5134
rect 59836 5070 59838 5122
rect 59890 5070 59892 5122
rect 59836 4564 59892 5070
rect 57372 4274 57428 4284
rect 59500 4452 59556 4462
rect 59500 4338 59556 4396
rect 59500 4286 59502 4338
rect 59554 4286 59556 4338
rect 59500 4274 59556 4286
rect 55468 4228 55524 4238
rect 55468 4134 55524 4172
rect 58380 4226 58436 4238
rect 58380 4174 58382 4226
rect 58434 4174 58436 4226
rect 54684 3666 54964 3668
rect 54684 3614 54686 3666
rect 54738 3614 54964 3666
rect 54684 3612 54964 3614
rect 54684 3602 54740 3612
rect 55468 3444 55524 3454
rect 55244 3388 55468 3444
rect 55244 800 55300 3388
rect 55468 3378 55524 3388
rect 55804 3444 55860 3454
rect 55804 3350 55860 3388
rect 56588 3444 56644 3454
rect 56588 3350 56644 3388
rect 57596 3444 57652 3454
rect 58156 3444 58212 3454
rect 57596 3442 58212 3444
rect 57596 3390 57598 3442
rect 57650 3390 58158 3442
rect 58210 3390 58212 3442
rect 57596 3388 58212 3390
rect 57596 3378 57652 3388
rect 57708 800 57764 3388
rect 58156 3378 58212 3388
rect 58380 800 58436 4174
rect 59500 3668 59556 3678
rect 59500 3574 59556 3612
rect 59836 800 59892 4508
rect 60060 4226 60116 32732
rect 60172 23828 60228 32956
rect 60396 32900 60452 41694
rect 60620 40964 60676 40974
rect 60956 40964 61012 41918
rect 60620 40962 61012 40964
rect 60620 40910 60622 40962
rect 60674 40910 61012 40962
rect 60620 40908 61012 40910
rect 60396 32834 60452 32844
rect 60508 40292 60564 40302
rect 60172 23762 60228 23772
rect 60060 4174 60062 4226
rect 60114 4174 60116 4226
rect 60060 4162 60116 4174
rect 60508 3668 60564 40236
rect 60620 38052 60676 40908
rect 61068 39060 61124 43260
rect 61180 41972 61236 43484
rect 61628 43484 61796 43540
rect 61852 44098 61908 44110
rect 61852 44046 61854 44098
rect 61906 44046 61908 44098
rect 61180 41906 61236 41916
rect 61292 43092 61348 43102
rect 61180 41300 61236 41310
rect 61180 40628 61236 41244
rect 61180 40514 61236 40572
rect 61180 40462 61182 40514
rect 61234 40462 61236 40514
rect 61180 40450 61236 40462
rect 61292 40290 61348 43036
rect 61516 42980 61572 42990
rect 61404 42644 61460 42654
rect 61404 42550 61460 42588
rect 61404 41300 61460 41310
rect 61404 41206 61460 41244
rect 61516 41298 61572 42924
rect 61628 42644 61684 43484
rect 61852 43428 61908 44046
rect 61964 43876 62020 44268
rect 61964 43538 62020 43820
rect 62188 43708 62244 44268
rect 62412 44324 62468 44334
rect 62412 44230 62468 44268
rect 61964 43486 61966 43538
rect 62018 43486 62020 43538
rect 61964 43474 62020 43486
rect 62076 43652 62244 43708
rect 62300 43764 62356 43774
rect 61628 42550 61684 42588
rect 61740 42866 61796 42878
rect 61740 42814 61742 42866
rect 61794 42814 61796 42866
rect 61740 42082 61796 42814
rect 61740 42030 61742 42082
rect 61794 42030 61796 42082
rect 61740 42018 61796 42030
rect 61852 42084 61908 43372
rect 62076 43316 62132 43652
rect 62300 43538 62356 43708
rect 62300 43486 62302 43538
rect 62354 43486 62356 43538
rect 62300 43474 62356 43486
rect 62412 43538 62468 43550
rect 62412 43486 62414 43538
rect 62466 43486 62468 43538
rect 62412 43316 62468 43486
rect 62076 43260 62244 43316
rect 62188 42866 62244 43260
rect 62412 43250 62468 43260
rect 62188 42814 62190 42866
rect 62242 42814 62244 42866
rect 62188 42802 62244 42814
rect 61852 42018 61908 42028
rect 61516 41246 61518 41298
rect 61570 41246 61572 41298
rect 61516 41234 61572 41246
rect 61628 40964 61684 40974
rect 62188 40964 62244 40974
rect 61628 40870 61684 40908
rect 61964 40962 62244 40964
rect 61964 40910 62190 40962
rect 62242 40910 62244 40962
rect 61964 40908 62244 40910
rect 61964 40628 62020 40908
rect 62188 40898 62244 40908
rect 61964 40534 62020 40572
rect 61516 40404 61572 40442
rect 61516 40338 61572 40348
rect 62412 40404 62468 40414
rect 62412 40310 62468 40348
rect 61292 40238 61294 40290
rect 61346 40238 61348 40290
rect 61292 40226 61348 40238
rect 62636 39396 62692 45164
rect 62748 44994 62804 45006
rect 62748 44942 62750 44994
rect 62802 44942 62804 44994
rect 62748 44548 62804 44942
rect 62748 44482 62804 44492
rect 62748 43540 62804 43550
rect 62748 43446 62804 43484
rect 62748 42868 62804 42878
rect 62860 42868 62916 45388
rect 62972 44882 63028 45948
rect 62972 44830 62974 44882
rect 63026 44830 63028 44882
rect 62972 44818 63028 44830
rect 63308 44548 63364 47406
rect 63532 46788 63588 50372
rect 63868 49026 63924 51324
rect 64092 51380 64148 52108
rect 64540 52098 64596 52108
rect 64876 51940 64932 55580
rect 65100 55412 65156 62132
rect 65324 61012 65380 62300
rect 65436 62290 65492 62300
rect 65548 62188 65604 63084
rect 65772 63138 65828 63150
rect 65772 63086 65774 63138
rect 65826 63086 65828 63138
rect 65772 62916 65828 63086
rect 66332 63028 66388 63038
rect 66444 63028 66500 64428
rect 66668 64594 66724 64606
rect 66668 64542 66670 64594
rect 66722 64542 66724 64594
rect 66556 64372 66612 64382
rect 66556 64146 66612 64316
rect 66556 64094 66558 64146
rect 66610 64094 66612 64146
rect 66556 64082 66612 64094
rect 66668 63812 66724 64542
rect 66668 63746 66724 63756
rect 66332 63026 66500 63028
rect 66332 62974 66334 63026
rect 66386 62974 66500 63026
rect 66332 62972 66500 62974
rect 66780 63252 66836 65548
rect 67116 64482 67172 66108
rect 67340 66050 67396 68012
rect 67788 67228 67844 113372
rect 68908 69188 68964 69198
rect 68908 67228 68964 69132
rect 69580 67228 69636 115388
rect 70140 115444 70196 115502
rect 70140 115378 70196 115388
rect 70700 90748 70756 115612
rect 71260 115556 71316 116396
rect 71372 116386 71428 116396
rect 72044 116340 72100 119200
rect 71708 115668 71764 115678
rect 71708 115574 71764 115612
rect 71148 115554 71316 115556
rect 71148 115502 71262 115554
rect 71314 115502 71316 115554
rect 71148 115500 71316 115502
rect 70700 90692 70868 90748
rect 67788 67172 68292 67228
rect 67340 65998 67342 66050
rect 67394 65998 67396 66050
rect 67340 64820 67396 65998
rect 67340 64754 67396 64764
rect 68012 64820 68068 64830
rect 68012 64726 68068 64764
rect 67676 64596 67732 64606
rect 67564 64594 67732 64596
rect 67564 64542 67678 64594
rect 67730 64542 67732 64594
rect 67564 64540 67732 64542
rect 67116 64430 67118 64482
rect 67170 64430 67172 64482
rect 67116 64036 67172 64430
rect 67116 63970 67172 63980
rect 67340 64484 67396 64494
rect 67340 64034 67396 64428
rect 67340 63982 67342 64034
rect 67394 63982 67396 64034
rect 66332 62962 66388 62972
rect 65772 62850 65828 62860
rect 65660 62356 65716 62366
rect 66780 62356 66836 63196
rect 67340 62580 67396 63982
rect 67564 63924 67620 64540
rect 67676 64530 67732 64540
rect 68124 64484 68180 64494
rect 67452 63812 67508 63822
rect 67452 63718 67508 63756
rect 67340 62514 67396 62524
rect 67564 62468 67620 63868
rect 67676 64148 67732 64158
rect 67676 63922 67732 64092
rect 68124 64146 68180 64428
rect 68124 64094 68126 64146
rect 68178 64094 68180 64146
rect 68124 64082 68180 64094
rect 67676 63870 67678 63922
rect 67730 63870 67732 63922
rect 67676 63858 67732 63870
rect 68012 63252 68068 63262
rect 68012 63158 68068 63196
rect 67564 62402 67620 62412
rect 65660 62262 65716 62300
rect 66556 62354 66836 62356
rect 66556 62302 66782 62354
rect 66834 62302 66836 62354
rect 66556 62300 66836 62302
rect 65548 62132 65828 62188
rect 65772 62130 65828 62132
rect 65772 62078 65774 62130
rect 65826 62078 65828 62130
rect 65772 61796 65828 62078
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65772 61740 66276 61796
rect 65212 60956 65380 61012
rect 65212 60676 65268 60956
rect 65660 60898 65716 60910
rect 65660 60846 65662 60898
rect 65714 60846 65716 60898
rect 65212 60610 65268 60620
rect 65324 60788 65380 60798
rect 65660 60788 65716 60846
rect 65380 60732 65716 60788
rect 65324 59106 65380 60732
rect 66220 60674 66276 61740
rect 66220 60622 66222 60674
rect 66274 60622 66276 60674
rect 65436 60564 65492 60574
rect 65436 60470 65492 60508
rect 65660 60564 65716 60574
rect 65324 59054 65326 59106
rect 65378 59054 65380 59106
rect 65324 58884 65380 59054
rect 65324 58818 65380 58828
rect 65548 59108 65604 59118
rect 65324 58658 65380 58670
rect 65324 58606 65326 58658
rect 65378 58606 65380 58658
rect 65324 58210 65380 58606
rect 65548 58324 65604 59052
rect 65548 58258 65604 58268
rect 65324 58158 65326 58210
rect 65378 58158 65380 58210
rect 65324 57876 65380 58158
rect 65324 57820 65604 57876
rect 65436 57540 65492 57550
rect 65324 57092 65380 57102
rect 65324 56998 65380 57036
rect 65436 56306 65492 57484
rect 65548 57204 65604 57820
rect 65548 57138 65604 57148
rect 65548 56980 65604 56990
rect 65548 56886 65604 56924
rect 65436 56254 65438 56306
rect 65490 56254 65492 56306
rect 65436 56242 65492 56254
rect 65548 56642 65604 56654
rect 65548 56590 65550 56642
rect 65602 56590 65604 56642
rect 65548 56532 65604 56590
rect 64988 55356 65156 55412
rect 65548 55636 65604 56476
rect 65548 55410 65604 55580
rect 65548 55358 65550 55410
rect 65602 55358 65604 55410
rect 64988 52388 65044 55356
rect 65548 55346 65604 55358
rect 65100 55188 65156 55198
rect 65100 55074 65156 55132
rect 65100 55022 65102 55074
rect 65154 55022 65156 55074
rect 65100 54292 65156 55022
rect 65100 54226 65156 54236
rect 65436 54402 65492 54414
rect 65436 54350 65438 54402
rect 65490 54350 65492 54402
rect 65436 53732 65492 54350
rect 65436 53666 65492 53676
rect 65660 53620 65716 60508
rect 65772 60562 65828 60574
rect 65772 60510 65774 60562
rect 65826 60510 65828 60562
rect 65772 60114 65828 60510
rect 66220 60562 66276 60622
rect 66220 60510 66222 60562
rect 66274 60510 66276 60562
rect 66220 60498 66276 60510
rect 66332 61348 66388 61358
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65772 60062 65774 60114
rect 65826 60062 65828 60114
rect 65772 60050 65828 60062
rect 66108 59332 66164 59342
rect 65772 59330 66164 59332
rect 65772 59278 66110 59330
rect 66162 59278 66164 59330
rect 65772 59276 66164 59278
rect 65772 58660 65828 59276
rect 66108 59266 66164 59276
rect 65884 59108 65940 59118
rect 65884 59014 65940 59052
rect 66220 59108 66276 59118
rect 66332 59108 66388 61292
rect 66220 59106 66388 59108
rect 66220 59054 66222 59106
rect 66274 59054 66388 59106
rect 66220 59052 66388 59054
rect 66556 60002 66612 62300
rect 66780 62290 66836 62300
rect 67452 62244 67508 62254
rect 67452 62242 67844 62244
rect 67452 62190 67454 62242
rect 67506 62190 67844 62242
rect 67452 62188 67844 62190
rect 67452 62178 67508 62188
rect 67788 62132 68180 62188
rect 67452 61908 67508 61918
rect 66668 61572 66724 61582
rect 66668 61478 66724 61516
rect 67228 61572 67284 61582
rect 66668 60676 66724 60686
rect 66668 60582 66724 60620
rect 66780 60564 66836 60574
rect 67228 60564 67284 61516
rect 67452 61570 67508 61852
rect 67452 61518 67454 61570
rect 67506 61518 67508 61570
rect 67452 61506 67508 61518
rect 67900 61684 67956 61694
rect 67900 61570 67956 61628
rect 67900 61518 67902 61570
rect 67954 61518 67956 61570
rect 67900 61506 67956 61518
rect 67564 61458 67620 61470
rect 67564 61406 67566 61458
rect 67618 61406 67620 61458
rect 67340 61348 67396 61358
rect 67340 61254 67396 61292
rect 67452 60900 67508 60910
rect 67564 60900 67620 61406
rect 67676 61348 67732 61358
rect 67676 61346 67956 61348
rect 67676 61294 67678 61346
rect 67730 61294 67956 61346
rect 67676 61292 67956 61294
rect 67676 61282 67732 61292
rect 67676 61124 67732 61134
rect 67676 61010 67732 61068
rect 67676 60958 67678 61010
rect 67730 60958 67732 61010
rect 67676 60946 67732 60958
rect 67452 60898 67620 60900
rect 67452 60846 67454 60898
rect 67506 60846 67620 60898
rect 67452 60844 67620 60846
rect 67452 60834 67508 60844
rect 67788 60786 67844 60798
rect 67788 60734 67790 60786
rect 67842 60734 67844 60786
rect 66780 60562 66948 60564
rect 66780 60510 66782 60562
rect 66834 60510 66948 60562
rect 66780 60508 66948 60510
rect 66780 60498 66836 60508
rect 66556 59950 66558 60002
rect 66610 59950 66612 60002
rect 66220 59042 66276 59052
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65772 58604 65940 58660
rect 65772 58324 65828 58334
rect 65772 58230 65828 58268
rect 65884 58212 65940 58604
rect 65884 58146 65940 58156
rect 66220 58212 66276 58222
rect 66220 58118 66276 58156
rect 65772 57652 65828 57662
rect 65772 57558 65828 57596
rect 66332 57652 66388 57662
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 66220 56980 66276 56990
rect 66332 56980 66388 57596
rect 66556 57652 66612 59950
rect 66780 60340 66836 60350
rect 66780 59442 66836 60284
rect 66780 59390 66782 59442
rect 66834 59390 66836 59442
rect 66780 59220 66836 59390
rect 66780 59154 66836 59164
rect 66556 57586 66612 57596
rect 66668 59108 66724 59118
rect 66220 56978 66388 56980
rect 66220 56926 66222 56978
rect 66274 56926 66388 56978
rect 66220 56924 66388 56926
rect 66444 57538 66500 57550
rect 66444 57486 66446 57538
rect 66498 57486 66500 57538
rect 66444 56980 66500 57486
rect 66220 56914 66276 56924
rect 66444 56914 66500 56924
rect 66668 57092 66724 59052
rect 66668 56754 66724 57036
rect 66892 56868 66948 60508
rect 67004 60452 67060 60462
rect 67004 60114 67060 60396
rect 67004 60062 67006 60114
rect 67058 60062 67060 60114
rect 67004 58884 67060 60062
rect 67228 60116 67284 60508
rect 67564 60676 67620 60686
rect 67452 60116 67508 60126
rect 67228 60114 67508 60116
rect 67228 60062 67454 60114
rect 67506 60062 67508 60114
rect 67228 60060 67508 60062
rect 67452 60050 67508 60060
rect 67564 59444 67620 60620
rect 67788 60228 67844 60734
rect 67900 60452 67956 61292
rect 68124 61124 68180 62132
rect 68124 61058 68180 61068
rect 68012 60900 68068 60910
rect 68012 60806 68068 60844
rect 67900 60386 67956 60396
rect 68012 60228 68068 60238
rect 67788 60226 68068 60228
rect 67788 60174 68014 60226
rect 68066 60174 68068 60226
rect 67788 60172 68068 60174
rect 68012 60162 68068 60172
rect 68124 59780 68180 59790
rect 68012 59778 68180 59780
rect 68012 59726 68126 59778
rect 68178 59726 68180 59778
rect 68012 59724 68180 59726
rect 67564 59442 67844 59444
rect 67564 59390 67566 59442
rect 67618 59390 67844 59442
rect 67564 59388 67844 59390
rect 67564 59378 67620 59388
rect 67116 59108 67172 59118
rect 67116 59014 67172 59052
rect 67004 58818 67060 58828
rect 67676 58996 67732 59006
rect 67564 58658 67620 58670
rect 67564 58606 67566 58658
rect 67618 58606 67620 58658
rect 67228 58436 67284 58446
rect 67228 58342 67284 58380
rect 67004 56980 67060 56990
rect 67004 56978 67396 56980
rect 67004 56926 67006 56978
rect 67058 56926 67396 56978
rect 67004 56924 67396 56926
rect 67004 56914 67060 56924
rect 66892 56802 66948 56812
rect 66668 56702 66670 56754
rect 66722 56702 66724 56754
rect 66332 56644 66388 56654
rect 65772 55972 65828 55982
rect 65772 55878 65828 55916
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65996 55412 66052 55422
rect 65996 55318 66052 55356
rect 66332 54740 66388 56588
rect 66668 56644 66724 56702
rect 67004 56756 67060 56766
rect 66668 56308 66724 56588
rect 66892 56644 66948 56654
rect 67004 56644 67060 56700
rect 66892 56642 67060 56644
rect 66892 56590 66894 56642
rect 66946 56590 67060 56642
rect 66892 56588 67060 56590
rect 66892 56578 66948 56588
rect 66668 56252 66948 56308
rect 66556 56082 66612 56094
rect 66556 56030 66558 56082
rect 66610 56030 66612 56082
rect 66556 55748 66612 56030
rect 66556 55682 66612 55692
rect 66668 56082 66724 56094
rect 66668 56030 66670 56082
rect 66722 56030 66724 56082
rect 66668 55412 66724 56030
rect 66668 55346 66724 55356
rect 66780 56082 66836 56094
rect 66780 56030 66782 56082
rect 66834 56030 66836 56082
rect 66332 54674 66388 54684
rect 66444 55076 66500 55086
rect 66780 55076 66836 56030
rect 66444 55074 66836 55076
rect 66444 55022 66446 55074
rect 66498 55022 66836 55074
rect 66444 55020 66836 55022
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65324 52834 65380 52846
rect 65324 52782 65326 52834
rect 65378 52782 65380 52834
rect 65324 52724 65380 52782
rect 64988 52322 65044 52332
rect 65212 52668 65380 52724
rect 65548 52834 65604 52846
rect 65548 52782 65550 52834
rect 65602 52782 65604 52834
rect 65100 52274 65156 52286
rect 65100 52222 65102 52274
rect 65154 52222 65156 52274
rect 64540 51884 64932 51940
rect 64988 52052 65044 52062
rect 64540 51490 64596 51884
rect 64540 51438 64542 51490
rect 64594 51438 64596 51490
rect 64540 51426 64596 51438
rect 64092 51378 64260 51380
rect 64092 51326 64094 51378
rect 64146 51326 64260 51378
rect 64092 51324 64260 51326
rect 64092 51314 64148 51324
rect 63980 51156 64036 51166
rect 63980 50820 64036 51100
rect 63980 50754 64036 50764
rect 64204 49924 64260 51324
rect 64764 51156 64820 51884
rect 64652 51100 64820 51156
rect 64876 51716 64932 51726
rect 64540 51044 64596 51054
rect 64428 50706 64484 50718
rect 64428 50654 64430 50706
rect 64482 50654 64484 50706
rect 64316 50484 64372 50522
rect 64316 50418 64372 50428
rect 64428 50034 64484 50654
rect 64540 50594 64596 50988
rect 64540 50542 64542 50594
rect 64594 50542 64596 50594
rect 64540 50530 64596 50542
rect 64428 49982 64430 50034
rect 64482 49982 64484 50034
rect 64428 49970 64484 49982
rect 64204 49830 64260 49868
rect 63980 49810 64036 49822
rect 63980 49758 63982 49810
rect 64034 49758 64036 49810
rect 63980 49140 64036 49758
rect 64092 49698 64148 49710
rect 64092 49646 64094 49698
rect 64146 49646 64148 49698
rect 64092 49364 64148 49646
rect 64652 49476 64708 51100
rect 64876 51044 64932 51660
rect 64876 50978 64932 50988
rect 64988 50596 65044 51996
rect 65100 51156 65156 52222
rect 65212 52162 65268 52668
rect 65212 52110 65214 52162
rect 65266 52110 65268 52162
rect 65212 51716 65268 52110
rect 65436 52052 65492 52062
rect 65436 51958 65492 51996
rect 65212 51650 65268 51660
rect 65436 51490 65492 51502
rect 65436 51438 65438 51490
rect 65490 51438 65492 51490
rect 65100 51090 65156 51100
rect 65212 51380 65268 51390
rect 64988 50530 65044 50540
rect 65100 50820 65156 50830
rect 64764 50372 64820 50382
rect 64764 50278 64820 50316
rect 64652 49420 64820 49476
rect 64092 49308 64708 49364
rect 63980 49074 64036 49084
rect 64652 49138 64708 49308
rect 64652 49086 64654 49138
rect 64706 49086 64708 49138
rect 64652 49074 64708 49086
rect 63868 48974 63870 49026
rect 63922 48974 63924 49026
rect 63868 48962 63924 48974
rect 64764 48692 64820 49420
rect 64428 48636 64820 48692
rect 64204 48468 64260 48478
rect 64204 48374 64260 48412
rect 63980 48244 64036 48254
rect 63980 48150 64036 48188
rect 64316 48242 64372 48254
rect 64316 48190 64318 48242
rect 64370 48190 64372 48242
rect 64316 48132 64372 48190
rect 64204 47684 64260 47694
rect 63532 46722 63588 46732
rect 63980 47572 64036 47582
rect 63980 47234 64036 47516
rect 63980 47182 63982 47234
rect 64034 47182 64036 47234
rect 63756 46676 63812 46686
rect 63756 46582 63812 46620
rect 63868 45780 63924 45790
rect 63868 45686 63924 45724
rect 63532 45332 63588 45342
rect 63308 44482 63364 44492
rect 63420 45106 63476 45118
rect 63420 45054 63422 45106
rect 63474 45054 63476 45106
rect 62972 44212 63028 44222
rect 62972 44118 63028 44156
rect 63420 44212 63476 45054
rect 63420 44146 63476 44156
rect 63196 44100 63252 44110
rect 63084 43652 63140 43662
rect 63084 43428 63140 43596
rect 63084 43362 63140 43372
rect 62748 42866 62916 42868
rect 62748 42814 62750 42866
rect 62802 42814 62916 42866
rect 62748 42812 62916 42814
rect 63196 42866 63252 44044
rect 63532 43764 63588 45276
rect 63980 44212 64036 47182
rect 64092 47348 64148 47358
rect 64092 46898 64148 47292
rect 64092 46846 64094 46898
rect 64146 46846 64148 46898
rect 64092 46834 64148 46846
rect 64092 46674 64148 46686
rect 64092 46622 64094 46674
rect 64146 46622 64148 46674
rect 64092 45892 64148 46622
rect 64092 45826 64148 45836
rect 64204 45330 64260 47628
rect 64316 47012 64372 48076
rect 64316 46946 64372 46956
rect 64204 45278 64206 45330
rect 64258 45278 64260 45330
rect 64204 45266 64260 45278
rect 64316 46676 64372 46686
rect 64428 46676 64484 48636
rect 64316 46674 64484 46676
rect 64316 46622 64318 46674
rect 64370 46622 64484 46674
rect 64316 46620 64484 46622
rect 64540 48468 64596 48478
rect 64316 45220 64372 46620
rect 64540 45332 64596 48412
rect 64540 45200 64596 45276
rect 64316 45154 64372 45164
rect 65100 44434 65156 50764
rect 65212 50706 65268 51324
rect 65212 50654 65214 50706
rect 65266 50654 65268 50706
rect 65212 50428 65268 50654
rect 65436 50708 65492 51438
rect 65436 50642 65492 50652
rect 65548 50428 65604 52782
rect 65660 51156 65716 53564
rect 66332 53956 66388 53966
rect 66220 53506 66276 53518
rect 66220 53454 66222 53506
rect 66274 53454 66276 53506
rect 66220 53396 66276 53454
rect 66220 53330 66276 53340
rect 66220 53172 66276 53182
rect 66332 53172 66388 53900
rect 66444 53508 66500 55020
rect 66892 54964 66948 56252
rect 66556 54908 66948 54964
rect 67116 56082 67172 56094
rect 67116 56030 67118 56082
rect 67170 56030 67172 56082
rect 66556 54628 66612 54908
rect 66556 54068 66612 54572
rect 67004 54628 67060 54638
rect 66556 54002 66612 54012
rect 66892 54516 66948 54526
rect 66892 53954 66948 54460
rect 66892 53902 66894 53954
rect 66946 53902 66948 53954
rect 66892 53890 66948 53902
rect 67004 53956 67060 54572
rect 67004 53824 67060 53900
rect 66444 53442 66500 53452
rect 66220 53170 66388 53172
rect 66220 53118 66222 53170
rect 66274 53118 66388 53170
rect 66220 53116 66388 53118
rect 67004 53284 67060 53294
rect 66220 53106 66276 53116
rect 65772 52946 65828 52958
rect 65772 52894 65774 52946
rect 65826 52894 65828 52946
rect 65772 52834 65828 52894
rect 66332 52948 66388 52958
rect 66332 52854 66388 52892
rect 66444 52946 66500 52958
rect 66444 52894 66446 52946
rect 66498 52894 66500 52946
rect 65772 52782 65774 52834
rect 65826 52782 65828 52834
rect 65772 52770 65828 52782
rect 66444 52836 66500 52894
rect 66892 52836 66948 52846
rect 66444 52834 66948 52836
rect 66444 52782 66894 52834
rect 66946 52782 66948 52834
rect 66444 52780 66948 52782
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65884 52388 65940 52398
rect 66444 52388 66500 52780
rect 66892 52770 66948 52780
rect 65772 51380 65828 51390
rect 65884 51380 65940 52332
rect 66332 52332 66500 52388
rect 66668 52388 66724 52398
rect 66220 51716 66276 51726
rect 66220 51602 66276 51660
rect 66220 51550 66222 51602
rect 66274 51550 66276 51602
rect 66220 51538 66276 51550
rect 65772 51378 65884 51380
rect 65772 51326 65774 51378
rect 65826 51326 65884 51378
rect 65772 51324 65884 51326
rect 65772 51314 65828 51324
rect 65884 51248 65940 51324
rect 65660 51100 65828 51156
rect 65660 50596 65716 50634
rect 65660 50530 65716 50540
rect 65212 50372 65380 50428
rect 65548 50372 65716 50428
rect 65324 50306 65380 50316
rect 65324 49700 65380 49710
rect 65324 49606 65380 49644
rect 65324 48692 65380 48702
rect 65324 46900 65380 48636
rect 65660 48468 65716 50372
rect 65772 49698 65828 51100
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65772 49646 65774 49698
rect 65826 49646 65828 49698
rect 65772 49252 65828 49646
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65772 49186 65828 49196
rect 65884 48468 65940 48478
rect 65660 48466 65940 48468
rect 65660 48414 65886 48466
rect 65938 48414 65940 48466
rect 65660 48412 65940 48414
rect 65884 48402 65940 48412
rect 66108 48242 66164 48254
rect 66108 48190 66110 48242
rect 66162 48190 66164 48242
rect 65100 44382 65102 44434
rect 65154 44382 65156 44434
rect 65100 44370 65156 44382
rect 65212 46898 65380 46900
rect 65212 46846 65326 46898
rect 65378 46846 65380 46898
rect 65212 46844 65380 46846
rect 63980 44146 64036 44156
rect 64204 44212 64260 44222
rect 63532 43650 63588 43708
rect 63532 43598 63534 43650
rect 63586 43598 63588 43650
rect 63532 43586 63588 43598
rect 63868 43876 63924 43886
rect 63196 42814 63198 42866
rect 63250 42814 63252 42866
rect 62748 42802 62804 42812
rect 63196 42802 63252 42814
rect 63532 42644 63588 42654
rect 63868 42644 63924 43820
rect 64204 43876 64260 44156
rect 64204 43810 64260 43820
rect 64540 43876 64596 43886
rect 64540 43762 64596 43820
rect 64540 43710 64542 43762
rect 64594 43710 64596 43762
rect 64540 43698 64596 43710
rect 63980 43426 64036 43438
rect 63980 43374 63982 43426
rect 64034 43374 64036 43426
rect 63980 42868 64036 43374
rect 63980 42802 64036 42812
rect 64428 43316 64484 43326
rect 64428 42866 64484 43260
rect 65212 43316 65268 46844
rect 65324 46834 65380 46844
rect 65548 48132 65604 48142
rect 65324 44994 65380 45006
rect 65324 44942 65326 44994
rect 65378 44942 65380 44994
rect 65324 44548 65380 44942
rect 65324 44482 65380 44492
rect 65324 43540 65380 43550
rect 65324 43446 65380 43484
rect 65212 43250 65268 43260
rect 64428 42814 64430 42866
rect 64482 42814 64484 42866
rect 64428 42802 64484 42814
rect 63980 42644 64036 42654
rect 63868 42642 64036 42644
rect 63868 42590 63982 42642
rect 64034 42590 64036 42642
rect 63868 42588 64036 42590
rect 63532 42550 63588 42588
rect 63980 42578 64036 42588
rect 63980 42194 64036 42206
rect 63980 42142 63982 42194
rect 64034 42142 64036 42194
rect 63980 42084 64036 42142
rect 63980 42018 64036 42028
rect 62748 40964 62804 40974
rect 62748 40870 62804 40908
rect 65548 39844 65604 48076
rect 65772 48020 65828 48030
rect 65772 47926 65828 47964
rect 66108 48020 66164 48190
rect 66108 47954 66164 47964
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 66332 47684 66388 52332
rect 66668 52162 66724 52332
rect 66668 52110 66670 52162
rect 66722 52110 66724 52162
rect 66556 51604 66612 51614
rect 66556 50594 66612 51548
rect 66556 50542 66558 50594
rect 66610 50542 66612 50594
rect 66556 50530 66612 50542
rect 66668 50428 66724 52110
rect 67004 52162 67060 53228
rect 67116 52276 67172 56030
rect 67340 55970 67396 56924
rect 67452 56644 67508 56654
rect 67452 56550 67508 56588
rect 67340 55918 67342 55970
rect 67394 55918 67396 55970
rect 67340 55906 67396 55918
rect 67340 55748 67396 55758
rect 67340 55410 67396 55692
rect 67340 55358 67342 55410
rect 67394 55358 67396 55410
rect 67340 55346 67396 55358
rect 67340 54404 67396 54414
rect 67452 54404 67508 54414
rect 67340 54402 67452 54404
rect 67340 54350 67342 54402
rect 67394 54350 67452 54402
rect 67340 54348 67452 54350
rect 67340 54338 67396 54348
rect 67340 54068 67396 54078
rect 67228 53730 67284 53742
rect 67228 53678 67230 53730
rect 67282 53678 67284 53730
rect 67228 52500 67284 53678
rect 67340 53730 67396 54012
rect 67340 53678 67342 53730
rect 67394 53678 67396 53730
rect 67340 53666 67396 53678
rect 67452 53732 67508 54348
rect 67228 52444 67396 52500
rect 67228 52276 67284 52286
rect 67116 52274 67284 52276
rect 67116 52222 67230 52274
rect 67282 52222 67284 52274
rect 67116 52220 67284 52222
rect 67228 52210 67284 52220
rect 67004 52110 67006 52162
rect 67058 52110 67060 52162
rect 66780 52052 66836 52062
rect 66780 51602 66836 51996
rect 66780 51550 66782 51602
rect 66834 51550 66836 51602
rect 66780 51538 66836 51550
rect 67004 51604 67060 52110
rect 67004 51538 67060 51548
rect 67228 51828 67284 51838
rect 67228 51602 67284 51772
rect 67228 51550 67230 51602
rect 67282 51550 67284 51602
rect 67228 51538 67284 51550
rect 67116 50820 67172 50830
rect 67116 50484 67172 50764
rect 67340 50818 67396 52444
rect 67452 52276 67508 53676
rect 67452 52210 67508 52220
rect 67564 52052 67620 58606
rect 67676 58546 67732 58940
rect 67676 58494 67678 58546
rect 67730 58494 67732 58546
rect 67676 58482 67732 58494
rect 67788 56532 67844 59388
rect 68012 59106 68068 59724
rect 68124 59714 68180 59724
rect 68012 59054 68014 59106
rect 68066 59054 68068 59106
rect 68012 57988 68068 59054
rect 68124 58658 68180 58670
rect 68124 58606 68126 58658
rect 68178 58606 68180 58658
rect 68124 58546 68180 58606
rect 68124 58494 68126 58546
rect 68178 58494 68180 58546
rect 68124 58482 68180 58494
rect 68012 57932 68180 57988
rect 67900 56868 67956 56878
rect 67900 56774 67956 56812
rect 67788 56466 67844 56476
rect 67788 56308 67844 56318
rect 67788 56306 67956 56308
rect 67788 56254 67790 56306
rect 67842 56254 67956 56306
rect 67788 56252 67956 56254
rect 67788 56242 67844 56252
rect 67788 55970 67844 55982
rect 67788 55918 67790 55970
rect 67842 55918 67844 55970
rect 67788 55860 67844 55918
rect 67788 55794 67844 55804
rect 67788 55522 67844 55534
rect 67788 55470 67790 55522
rect 67842 55470 67844 55522
rect 67788 55410 67844 55470
rect 67788 55358 67790 55410
rect 67842 55358 67844 55410
rect 67788 55346 67844 55358
rect 67900 54626 67956 56252
rect 68124 55412 68180 57932
rect 68236 56308 68292 67172
rect 68572 67172 68964 67228
rect 69468 67172 69636 67228
rect 68572 65378 68628 67172
rect 69244 66050 69300 66062
rect 69244 65998 69246 66050
rect 69298 65998 69300 66050
rect 68572 65326 68574 65378
rect 68626 65326 68628 65378
rect 68460 64708 68516 64718
rect 68460 64614 68516 64652
rect 68572 64148 68628 65326
rect 69132 65492 69188 65502
rect 69244 65492 69300 65998
rect 69132 65490 69300 65492
rect 69132 65438 69134 65490
rect 69186 65438 69300 65490
rect 69132 65436 69300 65438
rect 68684 64148 68740 64158
rect 68628 64146 68740 64148
rect 68628 64094 68686 64146
rect 68738 64094 68740 64146
rect 68628 64092 68740 64094
rect 68572 64016 68628 64092
rect 68684 64082 68740 64092
rect 69020 63810 69076 63822
rect 69020 63758 69022 63810
rect 69074 63758 69076 63810
rect 69020 63588 69076 63758
rect 69020 63522 69076 63532
rect 69132 63252 69188 65436
rect 69356 64708 69412 64718
rect 69356 64614 69412 64652
rect 69468 64148 69524 67172
rect 70252 66946 70308 66958
rect 70252 66894 70254 66946
rect 70306 66894 70308 66946
rect 70252 66836 70308 66894
rect 70252 66770 70308 66780
rect 70700 66946 70756 66958
rect 70700 66894 70702 66946
rect 70754 66894 70756 66946
rect 70700 66500 70756 66894
rect 70700 66434 70756 66444
rect 70476 66052 70532 66062
rect 69916 65380 69972 65390
rect 69580 65378 69972 65380
rect 69580 65326 69918 65378
rect 69970 65326 69972 65378
rect 69580 65324 69972 65326
rect 69580 64482 69636 65324
rect 69916 65314 69972 65324
rect 70476 64932 70532 65996
rect 70476 64866 70532 64876
rect 70700 65604 70756 65614
rect 69580 64430 69582 64482
rect 69634 64430 69636 64482
rect 69580 64418 69636 64430
rect 69692 64594 69748 64606
rect 69692 64542 69694 64594
rect 69746 64542 69748 64594
rect 69356 64092 69524 64148
rect 69356 63252 69412 64092
rect 69468 63924 69524 63934
rect 69692 63924 69748 64542
rect 69916 64596 69972 64606
rect 69916 64502 69972 64540
rect 70476 64594 70532 64606
rect 70476 64542 70478 64594
rect 70530 64542 70532 64594
rect 70476 64484 70532 64542
rect 70588 64596 70644 64606
rect 70588 64502 70644 64540
rect 70700 64594 70756 65548
rect 70700 64542 70702 64594
rect 70754 64542 70756 64594
rect 70700 64530 70756 64542
rect 70476 64418 70532 64428
rect 70700 64148 70756 64158
rect 70700 64054 70756 64092
rect 69524 63868 69748 63924
rect 70476 63924 70532 63934
rect 69468 63830 69524 63868
rect 70476 63830 70532 63868
rect 70140 63476 70196 63486
rect 69356 63196 69636 63252
rect 69132 63186 69188 63196
rect 68572 63028 68628 63038
rect 68460 62916 68516 62926
rect 68460 62822 68516 62860
rect 68572 62188 68628 62972
rect 69356 63028 69412 63038
rect 69356 62934 69412 62972
rect 69468 62916 69524 62926
rect 69468 62822 69524 62860
rect 69580 62244 69636 63196
rect 70140 63250 70196 63420
rect 70140 63198 70142 63250
rect 70194 63198 70196 63250
rect 70140 63028 70196 63198
rect 70140 62962 70196 62972
rect 68572 62132 68852 62188
rect 68348 61684 68404 61694
rect 68348 61590 68404 61628
rect 68572 61012 68628 61022
rect 68572 60918 68628 60956
rect 68684 60676 68740 60686
rect 68572 60674 68740 60676
rect 68572 60622 68686 60674
rect 68738 60622 68740 60674
rect 68572 60620 68740 60622
rect 68348 59778 68404 59790
rect 68348 59726 68350 59778
rect 68402 59726 68404 59778
rect 68348 59444 68404 59726
rect 68572 59556 68628 60620
rect 68684 60610 68740 60620
rect 68684 60452 68740 60462
rect 68684 60002 68740 60396
rect 68684 59950 68686 60002
rect 68738 59950 68740 60002
rect 68684 59938 68740 59950
rect 68572 59490 68628 59500
rect 68348 59378 68404 59388
rect 68460 59108 68516 59184
rect 68348 59052 68460 59108
rect 68348 58658 68404 59052
rect 68460 59042 68516 59052
rect 68572 58996 68628 59006
rect 68348 58606 68350 58658
rect 68402 58606 68404 58658
rect 68348 58594 68404 58606
rect 68460 58884 68516 58894
rect 68460 56868 68516 58828
rect 68572 58548 68628 58940
rect 68572 58416 68628 58492
rect 68572 57540 68628 57550
rect 68796 57540 68852 62132
rect 69580 62112 69636 62188
rect 70028 62580 70084 62590
rect 70028 61908 70084 62524
rect 70028 61842 70084 61852
rect 70476 62242 70532 62254
rect 70476 62190 70478 62242
rect 70530 62190 70532 62242
rect 70364 61684 70420 61694
rect 69468 61572 69524 61582
rect 69356 61570 69524 61572
rect 69356 61518 69470 61570
rect 69522 61518 69524 61570
rect 69356 61516 69524 61518
rect 69356 61012 69412 61516
rect 69468 61506 69524 61516
rect 69916 61572 69972 61582
rect 69916 61570 70308 61572
rect 69916 61518 69918 61570
rect 69970 61518 70308 61570
rect 69916 61516 70308 61518
rect 69916 61506 69972 61516
rect 70028 61348 70084 61358
rect 70028 61254 70084 61292
rect 70140 61346 70196 61358
rect 70140 61294 70142 61346
rect 70194 61294 70196 61346
rect 69356 60946 69412 60956
rect 69468 61010 69524 61022
rect 70140 61012 70196 61294
rect 69468 60958 69470 61010
rect 69522 60958 69524 61010
rect 69468 60564 69524 60958
rect 69580 60956 70196 61012
rect 69580 60786 69636 60956
rect 69580 60734 69582 60786
rect 69634 60734 69636 60786
rect 69580 60722 69636 60734
rect 69804 60788 69860 60798
rect 69804 60694 69860 60732
rect 69468 60498 69524 60508
rect 69356 60228 69412 60238
rect 69356 60002 69412 60172
rect 69916 60226 69972 60956
rect 70252 60900 70308 61516
rect 70252 60786 70308 60844
rect 70364 60898 70420 61628
rect 70364 60846 70366 60898
rect 70418 60846 70420 60898
rect 70364 60834 70420 60846
rect 70476 61012 70532 62190
rect 70252 60734 70254 60786
rect 70306 60734 70308 60786
rect 70252 60722 70308 60734
rect 69916 60174 69918 60226
rect 69970 60174 69972 60226
rect 69916 60162 69972 60174
rect 70364 60228 70420 60238
rect 69356 59950 69358 60002
rect 69410 59950 69412 60002
rect 69356 59938 69412 59950
rect 69580 60004 69636 60014
rect 69580 59778 69636 59948
rect 70028 59890 70084 59902
rect 70028 59838 70030 59890
rect 70082 59838 70084 59890
rect 69580 59726 69582 59778
rect 69634 59726 69636 59778
rect 68908 59556 68964 59566
rect 68908 59442 68964 59500
rect 68908 59390 68910 59442
rect 68962 59390 68964 59442
rect 68908 59378 68964 59390
rect 69356 59444 69412 59454
rect 69356 59350 69412 59388
rect 69468 59220 69524 59230
rect 69468 59126 69524 59164
rect 69356 59108 69412 59118
rect 69132 58884 69188 58894
rect 69132 57876 69188 58828
rect 69356 58546 69412 59052
rect 69580 58996 69636 59726
rect 69804 59778 69860 59790
rect 69804 59726 69806 59778
rect 69858 59726 69860 59778
rect 69692 59556 69748 59566
rect 69692 59442 69748 59500
rect 69692 59390 69694 59442
rect 69746 59390 69748 59442
rect 69692 59378 69748 59390
rect 69580 58930 69636 58940
rect 69804 58660 69860 59726
rect 70028 59780 70084 59838
rect 69916 59444 69972 59454
rect 69916 59350 69972 59388
rect 70028 59108 70084 59724
rect 70028 59042 70084 59052
rect 70140 59218 70196 59230
rect 70140 59166 70142 59218
rect 70194 59166 70196 59218
rect 69804 58594 69860 58604
rect 69916 58996 69972 59006
rect 69356 58494 69358 58546
rect 69410 58494 69412 58546
rect 69244 58436 69300 58446
rect 69356 58436 69412 58494
rect 69580 58548 69636 58558
rect 69300 58380 69412 58436
rect 69468 58436 69524 58446
rect 69244 58370 69300 58380
rect 69132 57820 69300 57876
rect 68572 57538 68852 57540
rect 68572 57486 68574 57538
rect 68626 57486 68852 57538
rect 68572 57484 68852 57486
rect 69132 57650 69188 57662
rect 69132 57598 69134 57650
rect 69186 57598 69188 57650
rect 68572 57474 68628 57484
rect 68460 56812 68740 56868
rect 68572 56642 68628 56654
rect 68572 56590 68574 56642
rect 68626 56590 68628 56642
rect 68572 56532 68628 56590
rect 68572 56466 68628 56476
rect 68460 56308 68516 56318
rect 68236 56306 68516 56308
rect 68236 56254 68462 56306
rect 68514 56254 68516 56306
rect 68236 56252 68516 56254
rect 68236 55522 68292 56252
rect 68460 56242 68516 56252
rect 68572 56308 68628 56318
rect 68572 56214 68628 56252
rect 68684 56306 68740 56812
rect 69132 56532 69188 57598
rect 69244 56978 69300 57820
rect 69468 57650 69524 58380
rect 69580 58434 69636 58492
rect 69580 58382 69582 58434
rect 69634 58382 69636 58434
rect 69580 58370 69636 58382
rect 69804 58324 69860 58334
rect 69916 58324 69972 58940
rect 70028 58884 70084 58894
rect 70028 58434 70084 58828
rect 70028 58382 70030 58434
rect 70082 58382 70084 58434
rect 70028 58370 70084 58382
rect 69804 58322 69972 58324
rect 69804 58270 69806 58322
rect 69858 58270 69972 58322
rect 69804 58268 69972 58270
rect 69804 58258 69860 58268
rect 70140 58212 70196 59166
rect 70364 59220 70420 60172
rect 70476 60114 70532 60956
rect 70476 60062 70478 60114
rect 70530 60062 70532 60114
rect 70476 60050 70532 60062
rect 70588 62244 70644 62254
rect 70588 59444 70644 62188
rect 70812 61908 70868 90692
rect 71148 64148 71204 115500
rect 71260 115490 71316 115500
rect 72044 114996 72100 116284
rect 72492 116562 72548 116574
rect 72492 116510 72494 116562
rect 72546 116510 72548 116562
rect 72380 115668 72436 115678
rect 72380 115574 72436 115612
rect 72156 114996 72212 115006
rect 72044 114994 72212 114996
rect 72044 114942 72158 114994
rect 72210 114942 72212 114994
rect 72044 114940 72212 114942
rect 72156 114930 72212 114940
rect 71260 94388 71316 94398
rect 71260 94294 71316 94332
rect 71820 94388 71876 94398
rect 71820 90748 71876 94332
rect 72156 94276 72212 94286
rect 72156 94182 72212 94220
rect 71820 90692 71988 90748
rect 71708 67732 71764 67742
rect 71372 67730 71764 67732
rect 71372 67678 71710 67730
rect 71762 67678 71764 67730
rect 71372 67676 71764 67678
rect 71372 67282 71428 67676
rect 71708 67666 71764 67676
rect 71372 67230 71374 67282
rect 71426 67230 71428 67282
rect 71372 67218 71428 67230
rect 71932 67228 71988 90692
rect 72380 68180 72436 68190
rect 71820 67172 71988 67228
rect 72044 67618 72100 67630
rect 72044 67566 72046 67618
rect 72098 67566 72100 67618
rect 71708 66834 71764 66846
rect 71708 66782 71710 66834
rect 71762 66782 71764 66834
rect 71708 66500 71764 66782
rect 71708 66434 71764 66444
rect 71372 66276 71428 66286
rect 71372 66274 71652 66276
rect 71372 66222 71374 66274
rect 71426 66222 71652 66274
rect 71372 66220 71652 66222
rect 71372 66210 71428 66220
rect 71260 64484 71316 64494
rect 71484 64484 71540 64494
rect 71316 64428 71428 64484
rect 71260 64352 71316 64428
rect 71148 64082 71204 64092
rect 71148 63924 71204 63934
rect 71204 63868 71316 63924
rect 71148 63830 71204 63868
rect 71036 62914 71092 62926
rect 71036 62862 71038 62914
rect 71090 62862 71092 62914
rect 71036 62356 71092 62862
rect 71148 62356 71204 62366
rect 71036 62300 71148 62356
rect 71148 62290 71204 62300
rect 70924 62244 70980 62254
rect 70980 62188 71092 62244
rect 70924 62150 70980 62188
rect 70812 61842 70868 61852
rect 70812 61684 70868 61694
rect 71036 61684 71092 62188
rect 70812 61682 71092 61684
rect 70812 61630 70814 61682
rect 70866 61630 71092 61682
rect 70812 61628 71092 61630
rect 71148 61684 71204 61694
rect 70812 61618 70868 61628
rect 71148 61572 71204 61628
rect 70924 61516 71204 61572
rect 70924 61458 70980 61516
rect 70924 61406 70926 61458
rect 70978 61406 70980 61458
rect 70924 61394 70980 61406
rect 70588 59378 70644 59388
rect 70700 61348 70756 61358
rect 70588 59220 70644 59230
rect 70364 59218 70644 59220
rect 70364 59166 70590 59218
rect 70642 59166 70644 59218
rect 70364 59164 70644 59166
rect 70364 58884 70420 59164
rect 70588 59154 70644 59164
rect 70364 58818 70420 58828
rect 70700 58434 70756 61292
rect 70924 60900 70980 60910
rect 70924 60806 70980 60844
rect 71036 60674 71092 60686
rect 71036 60622 71038 60674
rect 71090 60622 71092 60674
rect 71036 60004 71092 60622
rect 71260 60004 71316 63868
rect 71372 62356 71428 64428
rect 71372 60228 71428 62300
rect 71484 60788 71540 64428
rect 71596 63138 71652 66220
rect 71708 64484 71764 64494
rect 71708 64390 71764 64428
rect 71596 63086 71598 63138
rect 71650 63086 71652 63138
rect 71596 62188 71652 63086
rect 71708 62356 71764 62366
rect 71708 62262 71764 62300
rect 71596 62132 71764 62188
rect 71708 61570 71764 62132
rect 71708 61518 71710 61570
rect 71762 61518 71764 61570
rect 71708 61348 71764 61518
rect 71708 61282 71764 61292
rect 71596 60788 71652 60798
rect 71484 60786 71652 60788
rect 71484 60734 71598 60786
rect 71650 60734 71652 60786
rect 71484 60732 71652 60734
rect 71372 60172 71540 60228
rect 71372 60004 71428 60014
rect 71036 60002 71428 60004
rect 71036 59950 71374 60002
rect 71426 59950 71428 60002
rect 71036 59948 71428 59950
rect 70924 59780 70980 59790
rect 70924 59686 70980 59724
rect 70700 58382 70702 58434
rect 70754 58382 70756 58434
rect 70700 58370 70756 58382
rect 70812 59220 70868 59230
rect 70812 59108 70868 59164
rect 71036 59108 71092 59948
rect 71372 59938 71428 59948
rect 70812 59106 71092 59108
rect 70812 59054 71038 59106
rect 71090 59054 71092 59106
rect 70812 59052 71092 59054
rect 70364 58212 70420 58222
rect 70812 58212 70868 59052
rect 71036 59042 71092 59052
rect 71148 59780 71204 59790
rect 71484 59780 71540 60172
rect 70924 58546 70980 58558
rect 70924 58494 70926 58546
rect 70978 58494 70980 58546
rect 70924 58436 70980 58494
rect 70924 58370 70980 58380
rect 71036 58212 71092 58222
rect 70140 58210 70420 58212
rect 70140 58158 70366 58210
rect 70418 58158 70420 58210
rect 70140 58156 70420 58158
rect 69468 57598 69470 57650
rect 69522 57598 69524 57650
rect 69468 57586 69524 57598
rect 69692 57650 69748 57662
rect 69692 57598 69694 57650
rect 69746 57598 69748 57650
rect 69244 56926 69246 56978
rect 69298 56926 69300 56978
rect 69244 56914 69300 56926
rect 69580 57538 69636 57550
rect 69580 57486 69582 57538
rect 69634 57486 69636 57538
rect 69580 56980 69636 57486
rect 69580 56914 69636 56924
rect 69132 56466 69188 56476
rect 68684 56254 68686 56306
rect 68738 56254 68740 56306
rect 68348 56084 68404 56094
rect 68348 56082 68516 56084
rect 68348 56030 68350 56082
rect 68402 56030 68516 56082
rect 68348 56028 68516 56030
rect 68348 56018 68404 56028
rect 68460 55972 68516 56028
rect 68236 55470 68238 55522
rect 68290 55470 68292 55522
rect 68236 55458 68292 55470
rect 68348 55860 68404 55870
rect 68124 55346 68180 55356
rect 68236 55300 68292 55310
rect 68348 55300 68404 55804
rect 68236 55298 68404 55300
rect 68236 55246 68238 55298
rect 68290 55246 68404 55298
rect 68236 55244 68404 55246
rect 68236 55234 68292 55244
rect 67900 54574 67902 54626
rect 67954 54574 67956 54626
rect 67900 54562 67956 54574
rect 68012 54852 68068 54862
rect 68012 53844 68068 54796
rect 68460 54852 68516 55916
rect 68572 55412 68628 55422
rect 68684 55412 68740 56254
rect 69692 56308 69748 57598
rect 70252 57652 70308 57662
rect 70364 57652 70420 58156
rect 70700 58156 70868 58212
rect 70924 58210 71092 58212
rect 70924 58158 71038 58210
rect 71090 58158 71092 58210
rect 70924 58156 71092 58158
rect 70700 57762 70756 58156
rect 70812 57876 70868 57886
rect 70924 57876 70980 58156
rect 71036 58146 71092 58156
rect 71148 57988 71204 59724
rect 71372 59724 71540 59780
rect 71596 60116 71652 60732
rect 71820 60452 71876 67172
rect 72044 66386 72100 67566
rect 72380 67228 72436 68124
rect 72044 66334 72046 66386
rect 72098 66334 72100 66386
rect 72044 66322 72100 66334
rect 72156 67172 72212 67182
rect 72156 65604 72212 67116
rect 72268 67170 72324 67182
rect 72268 67118 72270 67170
rect 72322 67118 72324 67170
rect 72380 67162 72436 67172
rect 72268 67060 72324 67118
rect 72268 66994 72324 67004
rect 72380 67058 72436 67070
rect 72380 67006 72382 67058
rect 72434 67006 72436 67058
rect 72380 66836 72436 67006
rect 72380 66770 72436 66780
rect 72044 65380 72100 65390
rect 72156 65380 72212 65548
rect 72044 65378 72212 65380
rect 72044 65326 72046 65378
rect 72098 65326 72212 65378
rect 72044 65324 72212 65326
rect 72044 65314 72100 65324
rect 72156 64818 72212 65324
rect 72156 64766 72158 64818
rect 72210 64766 72212 64818
rect 72156 64754 72212 64766
rect 72380 63026 72436 63038
rect 72380 62974 72382 63026
rect 72434 62974 72436 63026
rect 72044 62580 72100 62590
rect 72380 62580 72436 62974
rect 72044 62578 72436 62580
rect 72044 62526 72046 62578
rect 72098 62526 72436 62578
rect 72044 62524 72436 62526
rect 72044 62514 72100 62524
rect 72044 62354 72100 62366
rect 72044 62302 72046 62354
rect 72098 62302 72100 62354
rect 72044 61684 72100 62302
rect 72380 62356 72436 62366
rect 72380 62262 72436 62300
rect 72044 61618 72100 61628
rect 72156 61908 72212 61918
rect 71932 61012 71988 61050
rect 71932 60946 71988 60956
rect 71932 60788 71988 60798
rect 71932 60694 71988 60732
rect 71820 60396 72100 60452
rect 71820 60116 71876 60126
rect 71596 60114 71876 60116
rect 71596 60062 71822 60114
rect 71874 60062 71876 60114
rect 71596 60060 71876 60062
rect 71260 58212 71316 58222
rect 71260 58118 71316 58156
rect 71372 58100 71428 59724
rect 71372 58034 71428 58044
rect 71484 59556 71540 59566
rect 71484 59106 71540 59500
rect 71484 59054 71486 59106
rect 71538 59054 71540 59106
rect 70812 57874 70980 57876
rect 70812 57822 70814 57874
rect 70866 57822 70980 57874
rect 70812 57820 70980 57822
rect 71036 57932 71204 57988
rect 70812 57810 70868 57820
rect 70700 57710 70702 57762
rect 70754 57710 70756 57762
rect 70252 57650 70420 57652
rect 70252 57598 70254 57650
rect 70306 57598 70420 57650
rect 70252 57596 70420 57598
rect 70252 57586 70308 57596
rect 70252 56866 70308 56878
rect 70252 56814 70254 56866
rect 70306 56814 70308 56866
rect 69692 56242 69748 56252
rect 70140 56308 70196 56318
rect 68908 56084 68964 56094
rect 68908 55990 68964 56028
rect 70140 56082 70196 56252
rect 70140 56030 70142 56082
rect 70194 56030 70196 56082
rect 70140 56018 70196 56030
rect 69580 55972 69636 55982
rect 69580 55970 69972 55972
rect 69580 55918 69582 55970
rect 69634 55918 69972 55970
rect 69580 55916 69972 55918
rect 69580 55906 69636 55916
rect 68572 55410 68740 55412
rect 68572 55358 68574 55410
rect 68626 55358 68740 55410
rect 68572 55356 68740 55358
rect 68572 55346 68628 55356
rect 68460 54786 68516 54796
rect 68684 55188 68740 55356
rect 69356 55524 69412 55534
rect 68684 54738 68740 55132
rect 68684 54686 68686 54738
rect 68738 54686 68740 54738
rect 68124 54626 68180 54638
rect 68124 54574 68126 54626
rect 68178 54574 68180 54626
rect 68124 54404 68180 54574
rect 68124 54338 68180 54348
rect 68236 54292 68292 54302
rect 68236 54290 68628 54292
rect 68236 54238 68238 54290
rect 68290 54238 68628 54290
rect 68236 54236 68628 54238
rect 68236 54226 68292 54236
rect 68124 53844 68180 53854
rect 68012 53842 68180 53844
rect 68012 53790 68126 53842
rect 68178 53790 68180 53842
rect 68012 53788 68180 53790
rect 68124 53778 68180 53788
rect 68012 53618 68068 53630
rect 68012 53566 68014 53618
rect 68066 53566 68068 53618
rect 68012 53172 68068 53566
rect 68236 53508 68292 53518
rect 68236 53414 68292 53452
rect 67900 53116 68012 53172
rect 67788 52948 67844 52958
rect 67340 50766 67342 50818
rect 67394 50766 67396 50818
rect 67340 50754 67396 50766
rect 67452 51996 67620 52052
rect 67676 52946 67844 52948
rect 67676 52894 67790 52946
rect 67842 52894 67844 52946
rect 67676 52892 67844 52894
rect 67676 52164 67732 52892
rect 67788 52882 67844 52892
rect 67788 52388 67844 52398
rect 67900 52388 67956 53116
rect 68012 53106 68068 53116
rect 68572 53058 68628 54236
rect 68572 53006 68574 53058
rect 68626 53006 68628 53058
rect 68572 52994 68628 53006
rect 68684 52836 68740 54686
rect 68908 55300 68964 55310
rect 68348 52780 68740 52836
rect 68796 54628 68852 54638
rect 67788 52386 68292 52388
rect 67788 52334 67790 52386
rect 67842 52334 68292 52386
rect 67788 52332 68292 52334
rect 67788 52322 67844 52332
rect 67228 50708 67284 50718
rect 67228 50614 67284 50652
rect 67116 50428 67396 50484
rect 66444 50370 66724 50428
rect 66444 50318 66670 50370
rect 66722 50318 66724 50370
rect 66444 50316 66724 50318
rect 66444 49812 66500 50316
rect 66668 50306 66724 50316
rect 66892 50370 66948 50382
rect 66892 50318 66894 50370
rect 66946 50318 66948 50370
rect 66444 48804 66500 49756
rect 66780 49810 66836 49822
rect 66780 49758 66782 49810
rect 66834 49758 66836 49810
rect 66780 49700 66836 49758
rect 66780 49634 66836 49644
rect 66892 49698 66948 50318
rect 66892 49646 66894 49698
rect 66946 49646 66948 49698
rect 66892 49634 66948 49646
rect 67228 49586 67284 49598
rect 67228 49534 67230 49586
rect 67282 49534 67284 49586
rect 66444 48738 66500 48748
rect 66780 49252 66836 49262
rect 66220 47348 66276 47358
rect 66332 47348 66388 47628
rect 66668 48132 66724 48142
rect 66668 47572 66724 48076
rect 66668 47506 66724 47516
rect 66444 47348 66500 47358
rect 66332 47292 66444 47348
rect 66220 47254 66276 47292
rect 66444 47282 66500 47292
rect 66668 47012 66724 47022
rect 65772 46900 65828 46910
rect 65772 46806 65828 46844
rect 66668 46898 66724 46956
rect 66668 46846 66670 46898
rect 66722 46846 66724 46898
rect 66668 46834 66724 46846
rect 66220 46788 66276 46798
rect 66220 46694 66276 46732
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65772 45220 65828 45230
rect 65772 45126 65828 45164
rect 66444 44994 66500 45006
rect 66444 44942 66446 44994
rect 66498 44942 66500 44994
rect 66444 44884 66500 44942
rect 66444 44818 66500 44828
rect 66780 44996 66836 49196
rect 66892 48802 66948 48814
rect 66892 48750 66894 48802
rect 66946 48750 66948 48802
rect 66892 48692 66948 48750
rect 66892 48626 66948 48636
rect 67116 48466 67172 48478
rect 67116 48414 67118 48466
rect 67170 48414 67172 48466
rect 67116 48356 67172 48414
rect 67116 48290 67172 48300
rect 67228 48354 67284 49534
rect 67228 48302 67230 48354
rect 67282 48302 67284 48354
rect 67228 48290 67284 48302
rect 67340 48242 67396 50428
rect 67452 49028 67508 51996
rect 67564 51604 67620 51614
rect 67564 51510 67620 51548
rect 67676 50372 67732 52108
rect 67900 51938 67956 51950
rect 67900 51886 67902 51938
rect 67954 51886 67956 51938
rect 67788 50596 67844 50606
rect 67788 50502 67844 50540
rect 67676 49140 67732 50316
rect 67900 49364 67956 51886
rect 68012 51938 68068 51950
rect 68012 51886 68014 51938
rect 68066 51886 68068 51938
rect 68012 51492 68068 51886
rect 68012 51426 68068 51436
rect 68124 51380 68180 51390
rect 68124 51286 68180 51324
rect 68236 50706 68292 52332
rect 68236 50654 68238 50706
rect 68290 50654 68292 50706
rect 68236 50642 68292 50654
rect 68124 49812 68180 49822
rect 68124 49718 68180 49756
rect 68348 49588 68404 52780
rect 68460 52276 68516 52286
rect 68460 50428 68516 52220
rect 68572 52276 68628 52286
rect 68796 52276 68852 54572
rect 68908 53844 68964 55244
rect 69356 54852 69412 55468
rect 69692 55412 69748 55422
rect 69692 55298 69748 55356
rect 69692 55246 69694 55298
rect 69746 55246 69748 55298
rect 69580 55188 69636 55198
rect 69580 55094 69636 55132
rect 69468 55076 69524 55086
rect 69468 54982 69524 55020
rect 69356 54796 69636 54852
rect 69132 54404 69188 54414
rect 68908 53778 68964 53788
rect 69020 54348 69132 54404
rect 68572 52274 68852 52276
rect 68572 52222 68574 52274
rect 68626 52222 68852 52274
rect 68572 52220 68852 52222
rect 68572 51828 68628 52220
rect 69020 52164 69076 54348
rect 69132 54272 69188 54348
rect 69244 53506 69300 53518
rect 69244 53454 69246 53506
rect 69298 53454 69300 53506
rect 69244 53172 69300 53454
rect 69244 53106 69300 53116
rect 68796 52108 69076 52164
rect 69244 52164 69300 52174
rect 68796 52052 68852 52108
rect 69244 52070 69300 52108
rect 68572 51762 68628 51772
rect 68684 51996 68852 52052
rect 68572 51604 68628 51614
rect 68572 50706 68628 51548
rect 68684 50820 68740 51996
rect 69468 51492 69524 51502
rect 69468 51398 69524 51436
rect 68908 51380 68964 51390
rect 68908 51286 68964 51324
rect 68684 50754 68740 50764
rect 68796 51154 68852 51166
rect 68796 51102 68798 51154
rect 68850 51102 68852 51154
rect 68796 50818 68852 51102
rect 68796 50766 68798 50818
rect 68850 50766 68852 50818
rect 68796 50754 68852 50766
rect 68572 50654 68574 50706
rect 68626 50654 68628 50706
rect 68572 50642 68628 50654
rect 69356 50594 69412 50606
rect 69356 50542 69358 50594
rect 69410 50542 69412 50594
rect 69356 50428 69412 50542
rect 68460 50372 68852 50428
rect 68572 50148 68628 50158
rect 68572 49700 68628 50092
rect 68572 49606 68628 49644
rect 67900 49308 68180 49364
rect 68012 49140 68068 49150
rect 67676 49138 68068 49140
rect 67676 49086 68014 49138
rect 68066 49086 68068 49138
rect 67676 49084 68068 49086
rect 68012 49074 68068 49084
rect 67452 48962 67508 48972
rect 67452 48804 67508 48842
rect 67452 48738 67508 48748
rect 67788 48804 67844 48814
rect 67340 48190 67342 48242
rect 67394 48190 67396 48242
rect 67004 48130 67060 48142
rect 67004 48078 67006 48130
rect 67058 48078 67060 48130
rect 67004 48020 67060 48078
rect 67004 47954 67060 47964
rect 67004 47458 67060 47470
rect 67004 47406 67006 47458
rect 67058 47406 67060 47458
rect 67004 45668 67060 47406
rect 67228 46564 67284 46574
rect 67228 46470 67284 46508
rect 67228 46004 67284 46014
rect 67340 46004 67396 48190
rect 67452 48580 67508 48590
rect 67452 46116 67508 48524
rect 67676 48468 67732 48478
rect 67788 48468 67844 48748
rect 67676 48466 67844 48468
rect 67676 48414 67678 48466
rect 67730 48414 67844 48466
rect 67676 48412 67844 48414
rect 67676 48402 67732 48412
rect 67900 48242 67956 48254
rect 67900 48190 67902 48242
rect 67954 48190 67956 48242
rect 67900 48132 67956 48190
rect 67900 48066 67956 48076
rect 67676 48020 67732 48030
rect 67676 47570 67732 47964
rect 67676 47518 67678 47570
rect 67730 47518 67732 47570
rect 67676 47506 67732 47518
rect 67564 47348 67620 47358
rect 67564 47254 67620 47292
rect 67788 47236 67844 47246
rect 67788 47142 67844 47180
rect 67452 46050 67508 46060
rect 68012 46676 68068 46686
rect 67228 46002 67396 46004
rect 67228 45950 67230 46002
rect 67282 45950 67396 46002
rect 67228 45948 67396 45950
rect 67228 45938 67284 45948
rect 68012 45780 68068 46620
rect 68012 45686 68068 45724
rect 67004 45602 67060 45612
rect 67564 45668 67620 45678
rect 66892 44996 66948 45006
rect 66780 44994 66948 44996
rect 66780 44942 66894 44994
rect 66946 44942 66948 44994
rect 66780 44940 66948 44942
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 66332 44660 66388 44670
rect 65660 44324 65716 44334
rect 65660 43764 65716 44268
rect 66108 44324 66164 44334
rect 66108 44230 66164 44268
rect 65660 43698 65716 43708
rect 66332 43876 66388 44604
rect 66220 43652 66276 43662
rect 66332 43652 66388 43820
rect 66220 43650 66388 43652
rect 66220 43598 66222 43650
rect 66274 43598 66388 43650
rect 66220 43596 66388 43598
rect 66668 44548 66724 44558
rect 66220 43586 66276 43596
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65548 39778 65604 39788
rect 61068 39058 62132 39060
rect 61068 39006 61070 39058
rect 61122 39006 62132 39058
rect 61068 39004 62132 39006
rect 61068 38994 61124 39004
rect 62076 38834 62132 39004
rect 62076 38782 62078 38834
rect 62130 38782 62132 38834
rect 62076 38770 62132 38782
rect 62636 38834 62692 39340
rect 62972 39620 63028 39630
rect 62860 38948 62916 38958
rect 62860 38854 62916 38892
rect 62636 38782 62638 38834
rect 62690 38782 62692 38834
rect 62636 38770 62692 38782
rect 61740 38612 61796 38622
rect 61628 38610 61796 38612
rect 61628 38558 61742 38610
rect 61794 38558 61796 38610
rect 61628 38556 61796 38558
rect 61404 38052 61460 38062
rect 60620 38050 61460 38052
rect 60620 37998 61406 38050
rect 61458 37998 61460 38050
rect 60620 37996 61460 37998
rect 60620 37826 60676 37996
rect 61404 37986 61460 37996
rect 60620 37774 60622 37826
rect 60674 37774 60676 37826
rect 60620 32004 60676 37774
rect 61628 37266 61684 38556
rect 61740 38546 61796 38556
rect 62188 37940 62244 37950
rect 61852 37938 62244 37940
rect 61852 37886 62190 37938
rect 62242 37886 62244 37938
rect 61852 37884 62244 37886
rect 61852 37490 61908 37884
rect 62188 37874 62244 37884
rect 61852 37438 61854 37490
rect 61906 37438 61908 37490
rect 61852 37426 61908 37438
rect 61628 37214 61630 37266
rect 61682 37214 61684 37266
rect 61628 37202 61684 37214
rect 60620 31938 60676 31948
rect 62748 26516 62804 26526
rect 62748 26290 62804 26460
rect 62748 26238 62750 26290
rect 62802 26238 62804 26290
rect 62748 26226 62804 26238
rect 62748 5124 62804 5134
rect 61068 4564 61124 4574
rect 61068 4450 61124 4508
rect 61068 4398 61070 4450
rect 61122 4398 61124 4450
rect 61068 4386 61124 4398
rect 60508 3602 60564 3612
rect 62748 3444 62804 5068
rect 62972 4562 63028 39564
rect 63420 39396 63476 39406
rect 63420 39058 63476 39340
rect 63420 39006 63422 39058
rect 63474 39006 63476 39058
rect 63420 38994 63476 39006
rect 63868 38948 63924 38958
rect 63868 38164 63924 38892
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 64316 38164 64372 38174
rect 63868 38162 64372 38164
rect 63868 38110 64318 38162
rect 64370 38110 64372 38162
rect 63868 38108 64372 38110
rect 64316 31948 64372 38108
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 66668 31948 66724 44492
rect 66780 42868 66836 44940
rect 66892 44930 66948 44940
rect 67228 44884 67284 44894
rect 66892 44324 66948 44334
rect 66892 44230 66948 44268
rect 67228 44322 67284 44828
rect 67228 44270 67230 44322
rect 67282 44270 67284 44322
rect 67228 44258 67284 44270
rect 67452 44210 67508 44222
rect 67452 44158 67454 44210
rect 67506 44158 67508 44210
rect 67004 44100 67060 44110
rect 67004 44006 67060 44044
rect 67116 44098 67172 44110
rect 67116 44046 67118 44098
rect 67170 44046 67172 44098
rect 67116 43988 67172 44046
rect 67116 43922 67172 43932
rect 67452 43764 67508 44158
rect 67452 43698 67508 43708
rect 66780 42802 66836 42812
rect 64316 31892 65380 31948
rect 66668 31892 66836 31948
rect 63196 26516 63252 26526
rect 63196 26422 63252 26460
rect 63868 23828 63924 23838
rect 63868 8372 63924 23772
rect 63868 8370 64484 8372
rect 63868 8318 63870 8370
rect 63922 8318 64484 8370
rect 63868 8316 64484 8318
rect 63868 8306 63924 8316
rect 64428 8258 64484 8316
rect 64428 8206 64430 8258
rect 64482 8206 64484 8258
rect 64428 8194 64484 8206
rect 64764 8036 64820 8046
rect 64764 7942 64820 7980
rect 63980 5124 64036 5134
rect 63980 5030 64036 5068
rect 62972 4510 62974 4562
rect 63026 4510 63028 4562
rect 62972 4340 63028 4510
rect 65324 4562 65380 31892
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65324 4510 65326 4562
rect 65378 4510 65380 4562
rect 63420 4340 63476 4350
rect 62972 4338 63476 4340
rect 62972 4286 63422 4338
rect 63474 4286 63476 4338
rect 62972 4284 63476 4286
rect 63420 4274 63476 4284
rect 64092 4226 64148 4238
rect 64092 4174 64094 4226
rect 64146 4174 64148 4226
rect 63868 3780 63924 3790
rect 63756 3724 63868 3780
rect 63756 3666 63812 3724
rect 63868 3714 63924 3724
rect 63756 3614 63758 3666
rect 63810 3614 63812 3666
rect 63756 3602 63812 3614
rect 62636 3442 62804 3444
rect 62636 3390 62750 3442
rect 62802 3390 62804 3442
rect 62636 3388 62804 3390
rect 62636 800 62692 3388
rect 62748 3378 62804 3388
rect 63308 3444 63364 3454
rect 63308 800 63364 3388
rect 64092 3444 64148 4174
rect 64988 3556 65044 3566
rect 65324 3556 65380 4510
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 66780 3780 66836 31892
rect 67564 30100 67620 45612
rect 67900 44436 67956 44446
rect 68124 44436 68180 49308
rect 68348 49138 68404 49532
rect 68348 49086 68350 49138
rect 68402 49086 68404 49138
rect 68348 48804 68404 49086
rect 68348 48738 68404 48748
rect 68460 48356 68516 48366
rect 68460 48262 68516 48300
rect 68796 48244 68852 50372
rect 68684 48130 68740 48142
rect 68684 48078 68686 48130
rect 68738 48078 68740 48130
rect 68348 47572 68404 47582
rect 68348 47478 68404 47516
rect 68684 46786 68740 48078
rect 68684 46734 68686 46786
rect 68738 46734 68740 46786
rect 68684 46722 68740 46734
rect 68796 45108 68852 48188
rect 69020 50372 69412 50428
rect 69580 50428 69636 54796
rect 69692 54404 69748 55246
rect 69916 55300 69972 55916
rect 70028 55300 70084 55310
rect 69916 55298 70084 55300
rect 69916 55246 70030 55298
rect 70082 55246 70084 55298
rect 69916 55244 70084 55246
rect 70028 55234 70084 55244
rect 69804 54516 69860 54526
rect 70252 54516 70308 56814
rect 70364 55970 70420 57596
rect 70364 55918 70366 55970
rect 70418 55918 70420 55970
rect 70364 55906 70420 55918
rect 70476 57650 70532 57662
rect 70476 57598 70478 57650
rect 70530 57598 70532 57650
rect 70476 57092 70532 57598
rect 70588 57092 70644 57102
rect 70476 57036 70588 57092
rect 70364 55300 70420 55338
rect 70364 55234 70420 55244
rect 69804 54514 70308 54516
rect 69804 54462 69806 54514
rect 69858 54462 70308 54514
rect 69804 54460 70308 54462
rect 69804 54450 69860 54460
rect 69692 54338 69748 54348
rect 70140 54292 70196 54302
rect 70140 53842 70196 54236
rect 70140 53790 70142 53842
rect 70194 53790 70196 53842
rect 70140 53778 70196 53790
rect 70028 53732 70084 53742
rect 70028 53638 70084 53676
rect 69692 52836 69748 52846
rect 69692 52388 69748 52780
rect 69692 52274 69748 52332
rect 69692 52222 69694 52274
rect 69746 52222 69748 52274
rect 69692 52210 69748 52222
rect 70252 52276 70308 54460
rect 70364 55074 70420 55086
rect 70364 55022 70366 55074
rect 70418 55022 70420 55074
rect 70364 53954 70420 55022
rect 70476 54628 70532 57036
rect 70588 57026 70644 57036
rect 70700 56308 70756 57710
rect 71036 57652 71092 57932
rect 71484 57876 71540 59054
rect 70700 56242 70756 56252
rect 70812 57596 71092 57652
rect 71260 57820 71540 57876
rect 70588 55300 70644 55310
rect 70588 55206 70644 55244
rect 70476 54572 70644 54628
rect 70476 54404 70532 54414
rect 70476 54310 70532 54348
rect 70588 54180 70644 54572
rect 70364 53902 70366 53954
rect 70418 53902 70420 53954
rect 70364 53890 70420 53902
rect 70476 54124 70644 54180
rect 70476 53732 70532 54124
rect 70252 52210 70308 52220
rect 70364 53676 70532 53732
rect 69916 51380 69972 51390
rect 69916 51266 69972 51324
rect 69916 51214 69918 51266
rect 69970 51214 69972 51266
rect 69916 50484 69972 51214
rect 69580 50372 69748 50428
rect 69916 50418 69972 50428
rect 70140 50482 70196 50494
rect 70140 50430 70142 50482
rect 70194 50430 70196 50482
rect 69020 49698 69076 50372
rect 69020 49646 69022 49698
rect 69074 49646 69076 49698
rect 69020 46676 69076 49646
rect 69580 49140 69636 49150
rect 69692 49140 69748 50372
rect 70028 50036 70084 50046
rect 70140 50036 70196 50430
rect 70364 50428 70420 53676
rect 70588 53060 70644 53070
rect 70476 51268 70532 51278
rect 70476 51174 70532 51212
rect 70028 50034 70196 50036
rect 70028 49982 70030 50034
rect 70082 49982 70196 50034
rect 70028 49980 70196 49982
rect 70252 50372 70420 50428
rect 70588 50428 70644 53004
rect 70700 52836 70756 52846
rect 70700 52742 70756 52780
rect 70700 52276 70756 52286
rect 70700 52162 70756 52220
rect 70700 52110 70702 52162
rect 70754 52110 70756 52162
rect 70700 52098 70756 52110
rect 70812 50428 70868 57596
rect 71148 57538 71204 57550
rect 71148 57486 71150 57538
rect 71202 57486 71204 57538
rect 70924 56980 70980 56990
rect 70924 56886 70980 56924
rect 71148 56308 71204 57486
rect 71260 57092 71316 57820
rect 71596 57764 71652 60060
rect 71820 60050 71876 60060
rect 72044 59668 72100 60396
rect 71820 59612 72100 59668
rect 71260 57026 71316 57036
rect 71372 57708 71652 57764
rect 71708 58212 71764 58222
rect 71148 56242 71204 56252
rect 71036 55972 71092 55982
rect 71036 55878 71092 55916
rect 71036 55188 71092 55198
rect 71036 55094 71092 55132
rect 71260 53732 71316 53742
rect 71260 53638 71316 53676
rect 70924 53508 70980 53518
rect 70924 53414 70980 53452
rect 71372 52948 71428 57708
rect 71596 57538 71652 57550
rect 71596 57486 71598 57538
rect 71650 57486 71652 57538
rect 71596 57092 71652 57486
rect 71596 57026 71652 57036
rect 71484 56084 71540 56094
rect 71484 55970 71540 56028
rect 71484 55918 71486 55970
rect 71538 55918 71540 55970
rect 71484 55524 71540 55918
rect 71484 55458 71540 55468
rect 71708 55412 71764 58156
rect 71708 55346 71764 55356
rect 71484 55300 71540 55310
rect 71484 55206 71540 55244
rect 70924 52892 71428 52948
rect 70924 51492 70980 52892
rect 71372 52052 71428 52062
rect 71148 52050 71428 52052
rect 71148 51998 71374 52050
rect 71426 51998 71428 52050
rect 71148 51996 71428 51998
rect 71148 51602 71204 51996
rect 71372 51986 71428 51996
rect 71148 51550 71150 51602
rect 71202 51550 71204 51602
rect 71148 51538 71204 51550
rect 70924 51490 71092 51492
rect 70924 51438 70926 51490
rect 70978 51438 71092 51490
rect 70924 51436 71092 51438
rect 70924 51426 70980 51436
rect 71036 50428 71092 51436
rect 71148 51378 71204 51390
rect 71148 51326 71150 51378
rect 71202 51326 71204 51378
rect 71148 51268 71204 51326
rect 71484 51380 71540 51390
rect 71484 51286 71540 51324
rect 71148 51202 71204 51212
rect 71820 50428 71876 59612
rect 72044 59444 72100 59454
rect 72044 59350 72100 59388
rect 72044 58100 72100 58110
rect 71932 56308 71988 56318
rect 71932 55972 71988 56252
rect 71932 55878 71988 55916
rect 71932 55076 71988 55086
rect 71932 54982 71988 55020
rect 72044 51604 72100 58044
rect 72156 52836 72212 61852
rect 72380 61458 72436 61470
rect 72380 61406 72382 61458
rect 72434 61406 72436 61458
rect 72380 61012 72436 61406
rect 72380 60946 72436 60956
rect 72268 60786 72324 60798
rect 72268 60734 72270 60786
rect 72322 60734 72324 60786
rect 72268 60676 72324 60734
rect 72268 60610 72324 60620
rect 72492 56868 72548 116510
rect 73388 115892 73444 119200
rect 75404 116564 75460 119200
rect 75404 116498 75460 116508
rect 76300 116452 76356 116462
rect 76188 116450 76356 116452
rect 76188 116398 76302 116450
rect 76354 116398 76356 116450
rect 76188 116396 76356 116398
rect 74396 116340 74452 116350
rect 74396 116246 74452 116284
rect 75516 116228 75572 116238
rect 75516 116134 75572 116172
rect 76188 116228 76244 116396
rect 76300 116386 76356 116396
rect 73388 115826 73444 115836
rect 74172 115892 74228 115902
rect 72604 115778 72660 115790
rect 72604 115726 72606 115778
rect 72658 115726 72660 115778
rect 72604 115668 72660 115726
rect 73500 115668 73556 115678
rect 72604 115666 73556 115668
rect 72604 115614 73502 115666
rect 73554 115614 73556 115666
rect 72604 115612 73556 115614
rect 73500 115602 73556 115612
rect 74172 115554 74228 115836
rect 74172 115502 74174 115554
rect 74226 115502 74228 115554
rect 74172 115490 74228 115502
rect 74732 113428 74788 113438
rect 73948 106260 74004 106270
rect 73948 103012 74004 106204
rect 73948 102946 74004 102956
rect 74732 93492 74788 113372
rect 74732 93426 74788 93436
rect 74732 87332 74788 87342
rect 73276 67060 73332 67070
rect 73276 66946 73332 67004
rect 73276 66894 73278 66946
rect 73330 66894 73332 66946
rect 73276 66500 73332 66894
rect 74284 67058 74340 67070
rect 74284 67006 74286 67058
rect 74338 67006 74340 67058
rect 74284 66948 74340 67006
rect 74284 66882 74340 66892
rect 74620 66836 74676 66846
rect 73276 66434 73332 66444
rect 74172 66500 74228 66510
rect 74172 66386 74228 66444
rect 74172 66334 74174 66386
rect 74226 66334 74228 66386
rect 74172 66322 74228 66334
rect 74620 66276 74676 66780
rect 74620 65490 74676 66220
rect 74732 65940 74788 87276
rect 76188 84978 76244 116172
rect 76748 115780 76804 119200
rect 76972 116564 77028 116574
rect 76972 116470 77028 116508
rect 78092 116564 78148 119200
rect 78092 116498 78148 116508
rect 78204 116450 78260 116462
rect 78204 116398 78206 116450
rect 78258 116398 78260 116450
rect 76748 115714 76804 115724
rect 77532 115780 77588 115790
rect 76860 115666 76916 115678
rect 76860 115614 76862 115666
rect 76914 115614 76916 115666
rect 76188 84926 76190 84978
rect 76242 84926 76244 84978
rect 75628 84868 75684 84878
rect 76188 84868 76244 84926
rect 75628 84866 76244 84868
rect 75628 84814 75630 84866
rect 75682 84814 76244 84866
rect 75628 84812 76244 84814
rect 75628 84802 75684 84812
rect 74844 67842 74900 67854
rect 74844 67790 74846 67842
rect 74898 67790 74900 67842
rect 74844 66498 74900 67790
rect 75068 67618 75124 67630
rect 75068 67566 75070 67618
rect 75122 67566 75124 67618
rect 74956 67172 75012 67182
rect 75068 67172 75124 67566
rect 76188 67228 76244 84812
rect 74956 67170 75124 67172
rect 74956 67118 74958 67170
rect 75010 67118 75124 67170
rect 74956 67116 75124 67118
rect 75852 67172 76244 67228
rect 76412 115556 76468 115566
rect 76860 115556 76916 115614
rect 76412 115554 76916 115556
rect 76412 115502 76414 115554
rect 76466 115502 76916 115554
rect 76412 115500 76916 115502
rect 77532 115554 77588 115724
rect 77532 115502 77534 115554
rect 77586 115502 77588 115554
rect 74956 67106 75012 67116
rect 74844 66446 74846 66498
rect 74898 66446 74900 66498
rect 74844 66434 74900 66446
rect 74956 66948 75012 66958
rect 74732 65874 74788 65884
rect 74620 65438 74622 65490
rect 74674 65438 74676 65490
rect 74620 65426 74676 65438
rect 74172 65380 74228 65390
rect 74172 64372 74228 65324
rect 74172 64306 74228 64316
rect 74956 65380 75012 66892
rect 75180 66274 75236 66286
rect 75180 66222 75182 66274
rect 75234 66222 75236 66274
rect 75068 65380 75124 65390
rect 74956 65378 75124 65380
rect 74956 65326 75070 65378
rect 75122 65326 75124 65378
rect 74956 65324 75124 65326
rect 73948 64260 74004 64270
rect 73388 63700 73444 63710
rect 73388 62468 73444 63644
rect 73388 60562 73444 62412
rect 73500 62356 73556 62366
rect 73500 62262 73556 62300
rect 73724 62356 73780 62366
rect 73724 62262 73780 62300
rect 73388 60510 73390 60562
rect 73442 60510 73444 60562
rect 73052 59780 73108 59790
rect 73388 59780 73444 60510
rect 73108 59724 73444 59780
rect 73500 61348 73556 61358
rect 73052 59686 73108 59724
rect 73052 57092 73108 57102
rect 73052 56978 73108 57036
rect 73052 56926 73054 56978
rect 73106 56926 73108 56978
rect 73052 56914 73108 56926
rect 72492 56802 72548 56812
rect 73500 56644 73556 61292
rect 73612 61012 73668 61022
rect 73612 60918 73668 60956
rect 73612 60676 73668 60686
rect 73612 60582 73668 60620
rect 73276 56642 73556 56644
rect 73276 56590 73502 56642
rect 73554 56590 73556 56642
rect 73276 56588 73556 56590
rect 72604 55972 72660 55982
rect 72604 54404 72660 55916
rect 72604 54310 72660 54348
rect 73276 54402 73332 56588
rect 73500 56578 73556 56588
rect 73276 54350 73278 54402
rect 73330 54350 73332 54402
rect 72156 52770 72212 52780
rect 73276 52276 73332 54350
rect 73276 52210 73332 52220
rect 73500 52274 73556 52286
rect 73500 52222 73502 52274
rect 73554 52222 73556 52274
rect 72044 51490 72100 51548
rect 73276 51604 73332 51614
rect 73276 51510 73332 51548
rect 72044 51438 72046 51490
rect 72098 51438 72100 51490
rect 70588 50372 70756 50428
rect 70812 50372 70980 50428
rect 71036 50372 71764 50428
rect 71820 50372 71988 50428
rect 70028 49970 70084 49980
rect 69804 49812 69860 49822
rect 69804 49718 69860 49756
rect 70028 49810 70084 49822
rect 70028 49758 70030 49810
rect 70082 49758 70084 49810
rect 70028 49140 70084 49758
rect 69580 49138 70084 49140
rect 69580 49086 69582 49138
rect 69634 49086 70084 49138
rect 69580 49084 70084 49086
rect 69580 49074 69636 49084
rect 69244 48692 69300 48702
rect 69244 48132 69300 48636
rect 70140 48244 70196 48254
rect 70140 48150 70196 48188
rect 69692 48132 69748 48142
rect 69244 48130 69412 48132
rect 69244 48078 69246 48130
rect 69298 48078 69412 48130
rect 69244 48076 69412 48078
rect 69244 48066 69300 48076
rect 69244 47348 69300 47358
rect 69244 47254 69300 47292
rect 69020 46610 69076 46620
rect 69356 46452 69412 48076
rect 69692 48038 69748 48076
rect 69804 47236 69860 47246
rect 69804 47142 69860 47180
rect 69356 46386 69412 46396
rect 68796 45042 68852 45052
rect 67900 44434 68180 44436
rect 67900 44382 67902 44434
rect 67954 44382 68180 44434
rect 67900 44380 68180 44382
rect 67900 44324 67956 44380
rect 67900 44258 67956 44268
rect 68460 44100 68516 44110
rect 68236 43764 68292 43774
rect 68236 43670 68292 43708
rect 68460 37828 68516 44044
rect 68460 37762 68516 37772
rect 67564 30034 67620 30044
rect 69356 30210 69412 30222
rect 69356 30158 69358 30210
rect 69410 30158 69412 30210
rect 69356 29988 69412 30158
rect 68124 28644 68180 28654
rect 68124 4564 68180 28588
rect 69356 26516 69412 29932
rect 70252 28644 70308 50372
rect 70364 49810 70420 49822
rect 70364 49758 70366 49810
rect 70418 49758 70420 49810
rect 70364 49700 70420 49758
rect 70364 49634 70420 49644
rect 70588 49250 70644 49262
rect 70588 49198 70590 49250
rect 70642 49198 70644 49250
rect 70588 49138 70644 49198
rect 70588 49086 70590 49138
rect 70642 49086 70644 49138
rect 70588 49074 70644 49086
rect 70588 48130 70644 48142
rect 70588 48078 70590 48130
rect 70642 48078 70644 48130
rect 70364 47460 70420 47470
rect 70588 47460 70644 48078
rect 70364 47458 70644 47460
rect 70364 47406 70366 47458
rect 70418 47406 70644 47458
rect 70364 47404 70644 47406
rect 70364 46676 70420 47404
rect 70364 46610 70420 46620
rect 70700 38668 70756 50372
rect 70812 50148 70868 50158
rect 70812 46562 70868 50092
rect 70924 49810 70980 50372
rect 70924 49758 70926 49810
rect 70978 49758 70980 49810
rect 70924 49250 70980 49758
rect 70924 49198 70926 49250
rect 70978 49198 70980 49250
rect 70924 49186 70980 49198
rect 71484 49812 71540 50372
rect 71708 50306 71764 50316
rect 71932 50148 71988 50372
rect 71932 50082 71988 50092
rect 72044 49924 72100 51438
rect 72156 51380 72212 51390
rect 72156 51286 72212 51324
rect 72380 51380 72436 51390
rect 72380 51286 72436 51324
rect 73500 51380 73556 52222
rect 73500 51268 73556 51324
rect 73724 51268 73780 51278
rect 73500 51266 73780 51268
rect 73500 51214 73726 51266
rect 73778 51214 73780 51266
rect 73500 51212 73780 51214
rect 73724 51156 73780 51212
rect 73724 51090 73780 51100
rect 72268 50708 72324 50718
rect 72268 50706 72548 50708
rect 72268 50654 72270 50706
rect 72322 50654 72548 50706
rect 72268 50652 72548 50654
rect 72268 50642 72324 50652
rect 72268 50484 72324 50494
rect 72268 50260 72324 50428
rect 72268 50204 72436 50260
rect 71484 49698 71540 49756
rect 71484 49646 71486 49698
rect 71538 49646 71540 49698
rect 71036 48804 71092 48814
rect 71148 48804 71204 48814
rect 71036 48802 71148 48804
rect 71036 48750 71038 48802
rect 71090 48750 71148 48802
rect 71036 48748 71148 48750
rect 71036 48738 71092 48748
rect 71148 47570 71204 48748
rect 71484 48804 71540 49646
rect 71820 49922 72100 49924
rect 71820 49870 72046 49922
rect 72098 49870 72100 49922
rect 71820 49868 72100 49870
rect 71820 49138 71876 49868
rect 72044 49858 72100 49868
rect 72268 49924 72324 49962
rect 72268 49858 72324 49868
rect 72268 49700 72324 49710
rect 72268 49606 72324 49644
rect 71820 49086 71822 49138
rect 71874 49086 71876 49138
rect 71820 49074 71876 49086
rect 71484 48738 71540 48748
rect 71148 47518 71150 47570
rect 71202 47518 71204 47570
rect 71148 47506 71204 47518
rect 70812 46510 70814 46562
rect 70866 46510 70868 46562
rect 70812 46498 70868 46510
rect 71372 45556 71428 45566
rect 70700 38612 70980 38668
rect 70252 28578 70308 28588
rect 69356 26450 69412 26460
rect 70812 26068 70868 26078
rect 69468 25844 69524 25854
rect 68796 22148 68852 22158
rect 68796 20580 68852 22092
rect 68796 20514 68852 20524
rect 68684 4564 68740 4574
rect 68124 4562 68740 4564
rect 68124 4510 68686 4562
rect 68738 4510 68740 4562
rect 68124 4508 68740 4510
rect 67788 4452 67844 4462
rect 67788 4358 67844 4396
rect 68124 4450 68180 4508
rect 68684 4498 68740 4508
rect 68124 4398 68126 4450
rect 68178 4398 68180 4450
rect 68124 4386 68180 4398
rect 66780 3714 66836 3724
rect 64988 3554 65380 3556
rect 64988 3502 64990 3554
rect 65042 3502 65380 3554
rect 64988 3500 65380 3502
rect 65436 3666 65492 3678
rect 65436 3614 65438 3666
rect 65490 3614 65492 3666
rect 64988 3490 65044 3500
rect 64092 3378 64148 3388
rect 64652 812 64820 868
rect 64652 800 64708 812
rect 43624 200 43848 728
rect 44968 200 45192 728
rect 46312 200 46536 728
rect 46620 700 46900 756
rect 46984 728 47236 800
rect 48328 728 48580 800
rect 49672 728 49924 800
rect 46984 200 47208 728
rect 48328 200 48552 728
rect 49672 200 49896 728
rect 50344 200 50568 800
rect 51688 728 51940 800
rect 51688 200 51912 728
rect 53032 200 53256 800
rect 54376 728 54628 800
rect 55048 728 55300 800
rect 54376 200 54600 728
rect 55048 200 55272 728
rect 56392 200 56616 800
rect 57708 728 57960 800
rect 58380 728 58632 800
rect 57736 200 57960 728
rect 58408 200 58632 728
rect 59752 200 59976 800
rect 61096 200 61320 800
rect 62440 728 62692 800
rect 63112 728 63364 800
rect 64456 728 64708 800
rect 64764 756 64820 812
rect 65436 756 65492 3614
rect 69468 3666 69524 25788
rect 70588 4452 70644 4462
rect 70364 4228 70420 4238
rect 70588 4228 70644 4396
rect 70364 4226 70644 4228
rect 70364 4174 70366 4226
rect 70418 4174 70644 4226
rect 70364 4172 70644 4174
rect 70364 4162 70420 4172
rect 69468 3614 69470 3666
rect 69522 3614 69524 3666
rect 69468 3602 69524 3614
rect 69020 3444 69076 3454
rect 69132 3444 69188 3454
rect 69020 3442 69132 3444
rect 69020 3390 69022 3442
rect 69074 3390 69132 3442
rect 69020 3388 69132 3390
rect 69020 3378 69076 3388
rect 69132 800 69188 3388
rect 70476 3444 70532 3454
rect 70476 3350 70532 3388
rect 70588 800 70644 4172
rect 70812 4226 70868 26012
rect 70924 25844 70980 38612
rect 71372 27748 71428 45500
rect 72268 30100 72324 30110
rect 72268 30006 72324 30044
rect 71372 27682 71428 27692
rect 72380 26068 72436 50204
rect 72492 49924 72548 50652
rect 72716 50594 72772 50606
rect 72716 50542 72718 50594
rect 72770 50542 72772 50594
rect 72716 50372 72772 50542
rect 72716 50306 72772 50316
rect 72492 49858 72548 49868
rect 73164 49924 73220 49934
rect 72380 26002 72436 26012
rect 73164 49700 73220 49868
rect 73276 49700 73332 49710
rect 73164 49698 73332 49700
rect 73164 49646 73278 49698
rect 73330 49646 73332 49698
rect 73164 49644 73332 49646
rect 70924 25778 70980 25788
rect 71820 4452 71876 4462
rect 71820 4358 71876 4396
rect 73164 4340 73220 49644
rect 73276 49634 73332 49644
rect 73724 48804 73780 48814
rect 73276 47572 73332 47582
rect 73276 46900 73332 47516
rect 73724 47570 73780 48748
rect 73724 47518 73726 47570
rect 73778 47518 73780 47570
rect 73724 47506 73780 47518
rect 73276 46834 73332 46844
rect 73948 43708 74004 64204
rect 74508 63250 74564 63262
rect 74508 63198 74510 63250
rect 74562 63198 74564 63250
rect 74172 62468 74228 62478
rect 74172 62374 74228 62412
rect 74508 62356 74564 63198
rect 74956 62914 75012 65324
rect 75068 65314 75124 65324
rect 75180 65380 75236 66222
rect 75628 66276 75684 66286
rect 75628 66182 75684 66220
rect 75180 65314 75236 65324
rect 75852 63476 75908 67172
rect 76300 66498 76356 66510
rect 76300 66446 76302 66498
rect 76354 66446 76356 66498
rect 75964 66164 76020 66174
rect 76300 66164 76356 66446
rect 75964 66162 76356 66164
rect 75964 66110 75966 66162
rect 76018 66110 76356 66162
rect 75964 66108 76356 66110
rect 75964 66098 76020 66108
rect 75852 63410 75908 63420
rect 74956 62862 74958 62914
rect 75010 62862 75012 62914
rect 74508 62290 74564 62300
rect 74732 62356 74788 62366
rect 74732 62262 74788 62300
rect 74508 61684 74564 61694
rect 74284 61628 74508 61684
rect 74172 61236 74228 61246
rect 74060 52276 74116 52286
rect 74060 52182 74116 52220
rect 73948 43652 74116 43708
rect 73948 43428 74004 43438
rect 73948 42868 74004 43372
rect 73948 42802 74004 42812
rect 74060 39620 74116 43652
rect 74060 39554 74116 39564
rect 73388 4340 73444 4350
rect 73164 4338 73444 4340
rect 73164 4286 73390 4338
rect 73442 4286 73444 4338
rect 73164 4284 73444 4286
rect 70812 4174 70814 4226
rect 70866 4174 70868 4226
rect 70812 4162 70868 4174
rect 72716 4228 72772 4238
rect 72716 800 72772 4172
rect 73164 3666 73220 4284
rect 73388 4274 73444 4284
rect 74060 4228 74116 4238
rect 74060 4134 74116 4172
rect 73164 3614 73166 3666
rect 73218 3614 73220 3666
rect 73164 3602 73220 3614
rect 74172 3666 74228 61180
rect 74284 61012 74340 61628
rect 74508 61590 74564 61628
rect 74956 61348 75012 62862
rect 74956 61254 75012 61292
rect 74284 60880 74340 60956
rect 76412 60004 76468 115500
rect 77532 115490 77588 115502
rect 78204 115220 78260 116398
rect 78764 115780 78820 119200
rect 78988 116564 79044 116574
rect 78988 116470 79044 116508
rect 79772 116564 79828 116574
rect 78764 115714 78820 115724
rect 78988 115780 79044 115790
rect 78988 115686 79044 115724
rect 77868 115164 78260 115220
rect 77868 114994 77924 115164
rect 77868 114942 77870 114994
rect 77922 114942 77924 114994
rect 76524 84868 76580 84878
rect 76524 84774 76580 84812
rect 77084 68852 77140 68862
rect 77084 66948 77140 68796
rect 77868 68852 77924 114942
rect 77868 68786 77924 68796
rect 77532 67842 77588 67854
rect 77532 67790 77534 67842
rect 77586 67790 77588 67842
rect 77532 67228 77588 67790
rect 77756 67788 78484 67844
rect 77756 67730 77812 67788
rect 77756 67678 77758 67730
rect 77810 67678 77812 67730
rect 77756 67666 77812 67678
rect 78316 67618 78372 67630
rect 78316 67566 78318 67618
rect 78370 67566 78372 67618
rect 77532 67172 77924 67228
rect 76524 66946 77140 66948
rect 76524 66894 77086 66946
rect 77138 66894 77140 66946
rect 76524 66892 77140 66894
rect 76524 66498 76580 66892
rect 77084 66882 77140 66892
rect 77644 67058 77700 67070
rect 77644 67006 77646 67058
rect 77698 67006 77700 67058
rect 77644 66948 77700 67006
rect 77644 66882 77700 66892
rect 76524 66446 76526 66498
rect 76578 66446 76580 66498
rect 76524 66386 76580 66446
rect 77868 66498 77924 67172
rect 78316 66948 78372 67566
rect 78428 67170 78484 67788
rect 78428 67118 78430 67170
rect 78482 67118 78484 67170
rect 78428 67106 78484 67118
rect 78316 66882 78372 66892
rect 77868 66446 77870 66498
rect 77922 66446 77924 66498
rect 77868 66434 77924 66446
rect 76524 66334 76526 66386
rect 76578 66334 76580 66386
rect 76524 66322 76580 66334
rect 78876 66388 78932 66398
rect 77420 66276 77476 66286
rect 77196 66164 77252 66174
rect 77196 66070 77252 66108
rect 77420 65714 77476 66220
rect 78204 66274 78260 66286
rect 78204 66222 78206 66274
rect 78258 66222 78260 66274
rect 78204 66164 78260 66222
rect 78204 66098 78260 66108
rect 78428 66276 78484 66286
rect 78428 66162 78484 66220
rect 78428 66110 78430 66162
rect 78482 66110 78484 66162
rect 77420 65662 77422 65714
rect 77474 65662 77476 65714
rect 77420 65650 77476 65662
rect 78428 65604 78484 66110
rect 78428 65538 78484 65548
rect 78652 66276 78708 66286
rect 76412 59938 76468 59948
rect 76636 60004 76692 60014
rect 76636 54628 76692 59948
rect 78652 56420 78708 66220
rect 78876 66162 78932 66332
rect 79548 66388 79604 66398
rect 79548 66294 79604 66332
rect 78876 66110 78878 66162
rect 78930 66110 78932 66162
rect 78876 66098 78932 66110
rect 78652 56354 78708 56364
rect 79772 56308 79828 116508
rect 81116 116564 81172 116574
rect 81228 116564 81284 119200
rect 81116 116562 81284 116564
rect 81116 116510 81118 116562
rect 81170 116510 81284 116562
rect 81116 116508 81284 116510
rect 81116 116498 81172 116508
rect 81228 116340 81284 116508
rect 81564 116564 81620 116574
rect 81564 116470 81620 116508
rect 81228 116274 81284 116284
rect 81276 116060 81540 116070
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81276 115994 81540 116004
rect 81788 115892 81844 115902
rect 81900 115892 81956 119200
rect 83468 116564 83524 119200
rect 84812 117012 84868 119200
rect 84812 116946 84868 116956
rect 83468 116498 83524 116508
rect 84812 116564 84868 116574
rect 84812 116470 84868 116508
rect 84140 116450 84196 116462
rect 84140 116398 84142 116450
rect 84194 116398 84196 116450
rect 82572 116340 82628 116350
rect 82572 116246 82628 116284
rect 81788 115890 81956 115892
rect 81788 115838 81790 115890
rect 81842 115838 81956 115890
rect 81788 115836 81956 115838
rect 81788 115826 81844 115836
rect 81900 115780 81956 115836
rect 81900 115714 81956 115724
rect 83244 115780 83300 115790
rect 83244 115686 83300 115724
rect 80108 115668 80164 115678
rect 80108 115666 80612 115668
rect 80108 115614 80110 115666
rect 80162 115614 80612 115666
rect 80108 115612 80612 115614
rect 80108 115602 80164 115612
rect 80556 115554 80612 115612
rect 80556 115502 80558 115554
rect 80610 115502 80612 115554
rect 80444 66948 80500 66958
rect 80444 61682 80500 66892
rect 80556 66946 80612 115502
rect 82236 115554 82292 115566
rect 82236 115502 82238 115554
rect 82290 115502 82292 115554
rect 81276 114492 81540 114502
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81276 114426 81540 114436
rect 81276 112924 81540 112934
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81276 112858 81540 112868
rect 81276 111356 81540 111366
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81276 111290 81540 111300
rect 81276 109788 81540 109798
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81276 109722 81540 109732
rect 81276 108220 81540 108230
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81276 108154 81540 108164
rect 81276 106652 81540 106662
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81276 106586 81540 106596
rect 81276 105084 81540 105094
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81276 105018 81540 105028
rect 81276 103516 81540 103526
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81276 103450 81540 103460
rect 81276 101948 81540 101958
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81276 101882 81540 101892
rect 81276 100380 81540 100390
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81276 100314 81540 100324
rect 81276 98812 81540 98822
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81276 98746 81540 98756
rect 81276 97244 81540 97254
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81276 97178 81540 97188
rect 81276 95676 81540 95686
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81276 95610 81540 95620
rect 81276 94108 81540 94118
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81276 94042 81540 94052
rect 81276 92540 81540 92550
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81276 92474 81540 92484
rect 81276 90972 81540 90982
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81276 90906 81540 90916
rect 81276 89404 81540 89414
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81276 89338 81540 89348
rect 81276 87836 81540 87846
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81276 87770 81540 87780
rect 81276 86268 81540 86278
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81276 86202 81540 86212
rect 81276 84700 81540 84710
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81276 84634 81540 84644
rect 81276 83132 81540 83142
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81276 83066 81540 83076
rect 81276 81564 81540 81574
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81276 81498 81540 81508
rect 81276 79996 81540 80006
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81276 79930 81540 79940
rect 81276 78428 81540 78438
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81276 78362 81540 78372
rect 81276 76860 81540 76870
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81276 76794 81540 76804
rect 81276 75292 81540 75302
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81276 75226 81540 75236
rect 81276 73724 81540 73734
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81276 73658 81540 73668
rect 81276 72156 81540 72166
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81276 72090 81540 72100
rect 81276 70588 81540 70598
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81276 70522 81540 70532
rect 81276 69020 81540 69030
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81276 68954 81540 68964
rect 81276 67452 81540 67462
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81276 67386 81540 67396
rect 82012 67058 82068 67070
rect 82012 67006 82014 67058
rect 82066 67006 82068 67058
rect 80556 66894 80558 66946
rect 80610 66894 80612 66946
rect 80556 66388 80612 66894
rect 81228 66948 81284 66958
rect 81228 66854 81284 66892
rect 80556 66322 80612 66332
rect 81676 66052 81732 66062
rect 81676 65958 81732 65996
rect 82012 66052 82068 67006
rect 82236 66276 82292 115502
rect 84140 115554 84196 116398
rect 84140 115502 84142 115554
rect 84194 115502 84196 115554
rect 83132 99876 83188 99886
rect 83132 68068 83188 99820
rect 83132 68002 83188 68012
rect 83244 79380 83300 79390
rect 82348 67284 82404 67322
rect 82348 67218 82404 67228
rect 82236 66210 82292 66220
rect 82012 65986 82068 65996
rect 81276 65884 81540 65894
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81276 65818 81540 65828
rect 81276 64316 81540 64326
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81276 64250 81540 64260
rect 81276 62748 81540 62758
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81276 62682 81540 62692
rect 80444 61630 80446 61682
rect 80498 61630 80500 61682
rect 80444 61618 80500 61630
rect 81116 61572 81172 61582
rect 81116 61478 81172 61516
rect 83020 61572 83076 61582
rect 83020 61478 83076 61516
rect 83244 61460 83300 79324
rect 83356 68068 83412 68078
rect 83356 66500 83412 68012
rect 83356 66434 83412 66444
rect 84140 61684 84196 115502
rect 85260 116452 85316 116462
rect 85260 115890 85316 116396
rect 85932 116452 85988 116462
rect 85932 116358 85988 116396
rect 85260 115838 85262 115890
rect 85314 115838 85316 115890
rect 85260 113428 85316 115838
rect 86156 115892 86212 119200
rect 86604 117012 86660 117022
rect 86604 116562 86660 116956
rect 86604 116510 86606 116562
rect 86658 116510 86660 116562
rect 86604 116498 86660 116510
rect 86156 115826 86212 115836
rect 86268 115666 86324 115678
rect 86268 115614 86270 115666
rect 86322 115614 86324 115666
rect 85820 115556 85876 115566
rect 86268 115556 86324 115614
rect 85820 115554 86324 115556
rect 85820 115502 85822 115554
rect 85874 115502 86324 115554
rect 85820 115500 86324 115502
rect 85820 115490 85876 115500
rect 85260 113362 85316 113372
rect 86268 68180 86324 115500
rect 86828 114772 86884 119200
rect 88172 116564 88228 119200
rect 88172 116498 88228 116508
rect 89068 116564 89124 116574
rect 89068 116470 89124 116508
rect 90860 116564 90916 119200
rect 90860 116498 90916 116508
rect 92652 116564 92708 116574
rect 92652 116470 92708 116508
rect 88284 116450 88340 116462
rect 88284 116398 88286 116450
rect 88338 116398 88340 116450
rect 86940 115892 86996 115902
rect 86940 115554 86996 115836
rect 87948 115668 88004 115678
rect 87948 115574 88004 115612
rect 88284 115668 88340 116398
rect 88284 115602 88340 115612
rect 89852 116452 89908 116462
rect 86940 115502 86942 115554
rect 86994 115502 86996 115554
rect 86940 115490 86996 115502
rect 86940 114772 86996 114782
rect 86828 114770 86996 114772
rect 86828 114718 86942 114770
rect 86994 114718 86996 114770
rect 86828 114716 86996 114718
rect 86940 114706 86996 114716
rect 88172 94612 88228 94622
rect 86268 68114 86324 68124
rect 86492 75684 86548 75694
rect 84140 61618 84196 61628
rect 83244 61394 83300 61404
rect 81276 61180 81540 61190
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81276 61114 81540 61124
rect 81276 59612 81540 59622
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81276 59546 81540 59556
rect 86492 58772 86548 75628
rect 86492 58706 86548 58716
rect 81276 58044 81540 58054
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81276 57978 81540 57988
rect 83132 57876 83188 57886
rect 79772 56242 79828 56252
rect 80108 56980 80164 56990
rect 76636 54562 76692 54572
rect 79436 56084 79492 56094
rect 79996 56084 80052 56094
rect 79436 56082 80052 56084
rect 79436 56030 79438 56082
rect 79490 56030 79998 56082
rect 80050 56030 80052 56082
rect 79436 56028 80052 56030
rect 79436 54516 79492 56028
rect 79996 56018 80052 56028
rect 79436 54450 79492 54460
rect 77868 53396 77924 53406
rect 76972 50708 77028 50718
rect 76972 48804 77028 50652
rect 75068 43428 75124 43438
rect 75068 29988 75124 43372
rect 75068 29894 75124 29932
rect 76524 30100 76580 30110
rect 76524 22482 76580 30044
rect 76524 22430 76526 22482
rect 76578 22430 76580 22482
rect 76524 22372 76580 22430
rect 76524 22306 76580 22316
rect 76524 4564 76580 4574
rect 76972 4564 77028 48748
rect 77868 24162 77924 53340
rect 79772 44436 79828 44446
rect 79772 24948 79828 44380
rect 80108 26292 80164 56924
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 80332 56196 80388 56206
rect 80332 56102 80388 56140
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 80556 48132 80612 48142
rect 80556 44884 80612 48076
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 80556 44818 80612 44828
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 82348 43428 82404 43438
rect 82348 43334 82404 43372
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 80108 26226 80164 26236
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 79772 24882 79828 24892
rect 77868 24110 77870 24162
rect 77922 24110 77924 24162
rect 77868 24050 77924 24110
rect 78428 24164 78484 24174
rect 78428 24162 78932 24164
rect 78428 24110 78430 24162
rect 78482 24110 78932 24162
rect 78428 24108 78932 24110
rect 78428 24098 78484 24108
rect 77868 23998 77870 24050
rect 77922 23998 77924 24050
rect 77868 23986 77924 23998
rect 78316 23716 78372 23726
rect 78316 23622 78372 23660
rect 77868 23266 77924 23278
rect 77868 23214 77870 23266
rect 77922 23214 77924 23266
rect 77644 23156 77700 23166
rect 77644 23062 77700 23100
rect 77868 22708 77924 23214
rect 78540 23156 78596 23166
rect 78540 23062 78596 23100
rect 78876 23154 78932 24108
rect 79100 23716 79156 23726
rect 79100 23266 79156 23660
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 79100 23214 79102 23266
rect 79154 23214 79156 23266
rect 79100 23202 79156 23214
rect 79660 23268 79716 23278
rect 79660 23266 80276 23268
rect 79660 23214 79662 23266
rect 79714 23214 80276 23266
rect 79660 23212 80276 23214
rect 79660 23202 79716 23212
rect 78876 23102 78878 23154
rect 78930 23102 78932 23154
rect 77868 22652 78372 22708
rect 78316 22482 78372 22652
rect 78316 22430 78318 22482
rect 78370 22430 78372 22482
rect 78316 22418 78372 22430
rect 77532 22372 77588 22382
rect 77532 21476 77588 22316
rect 77532 21410 77588 21420
rect 78876 8428 78932 23102
rect 80220 23042 80276 23212
rect 80220 22990 80222 23042
rect 80274 22990 80276 23042
rect 80220 22484 80276 22990
rect 80444 22484 80500 22494
rect 80220 22482 80612 22484
rect 80220 22430 80446 22482
rect 80498 22430 80612 22482
rect 80220 22428 80612 22430
rect 80444 22418 80500 22428
rect 76524 4562 77028 4564
rect 76524 4510 76526 4562
rect 76578 4510 77028 4562
rect 76524 4508 77028 4510
rect 76524 4498 76580 4508
rect 76972 4450 77028 4508
rect 78316 8372 78932 8428
rect 78316 4562 78372 8372
rect 78316 4510 78318 4562
rect 78370 4510 78372 4562
rect 76972 4398 76974 4450
rect 77026 4398 77028 4450
rect 76972 4386 77028 4398
rect 77308 4450 77364 4462
rect 77308 4398 77310 4450
rect 77362 4398 77364 4450
rect 74172 3614 74174 3666
rect 74226 3614 74228 3666
rect 74172 3602 74228 3614
rect 75740 4226 75796 4238
rect 75740 4174 75742 4226
rect 75794 4174 75796 4226
rect 74060 3444 74116 3454
rect 74060 800 74116 3388
rect 75068 3444 75124 3454
rect 75068 3350 75124 3388
rect 75740 3444 75796 4174
rect 77308 3556 77364 4398
rect 78316 4340 78372 4510
rect 80556 4562 80612 22428
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 83132 5908 83188 57820
rect 88172 55748 88228 94556
rect 88172 55682 88228 55692
rect 88508 58436 88564 58446
rect 88508 54516 88564 58380
rect 89852 57540 89908 116396
rect 91980 116450 92036 116462
rect 91980 116398 91982 116450
rect 92034 116398 92036 116450
rect 91196 116228 91252 116238
rect 91980 116228 92036 116398
rect 94220 116340 94276 119200
rect 94892 117348 94948 119200
rect 97580 117796 97636 119200
rect 97580 117740 97972 117796
rect 94892 117292 95172 117348
rect 95116 116562 95172 117292
rect 96636 116844 96900 116854
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96636 116778 96900 116788
rect 95116 116510 95118 116562
rect 95170 116510 95172 116562
rect 94332 116340 94388 116350
rect 94220 116338 94388 116340
rect 94220 116286 94334 116338
rect 94386 116286 94388 116338
rect 94220 116284 94388 116286
rect 94332 116274 94388 116284
rect 95116 116340 95172 116510
rect 95900 116562 95956 116574
rect 95900 116510 95902 116562
rect 95954 116510 95956 116562
rect 95900 116452 95956 116510
rect 95900 116386 95956 116396
rect 95116 116274 95172 116284
rect 96908 116340 96964 116350
rect 96908 116246 96964 116284
rect 97916 116338 97972 117740
rect 99148 116564 99204 116574
rect 99372 116564 99428 119200
rect 99148 116562 99428 116564
rect 99148 116510 99150 116562
rect 99202 116510 99428 116562
rect 99148 116508 99428 116510
rect 99148 116498 99204 116508
rect 97916 116286 97918 116338
rect 97970 116286 97972 116338
rect 97916 116274 97972 116286
rect 99372 116340 99428 116508
rect 99372 116274 99428 116284
rect 99820 116562 99876 116574
rect 99820 116510 99822 116562
rect 99874 116510 99876 116562
rect 91196 116226 92036 116228
rect 91196 116174 91198 116226
rect 91250 116174 92036 116226
rect 91196 116172 92036 116174
rect 91196 68068 91252 116172
rect 96636 115276 96900 115286
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96636 115210 96900 115220
rect 96636 113708 96900 113718
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96636 113642 96900 113652
rect 96636 112140 96900 112150
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96636 112074 96900 112084
rect 96636 110572 96900 110582
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96636 110506 96900 110516
rect 91196 68002 91252 68012
rect 93212 109284 93268 109294
rect 89852 57474 89908 57484
rect 91532 64708 91588 64718
rect 89964 54628 90020 54638
rect 89964 54534 90020 54572
rect 84812 54404 84868 54414
rect 83132 5842 83188 5852
rect 84140 27748 84196 27758
rect 81676 4900 81732 4910
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 80556 4510 80558 4562
rect 80610 4510 80612 4562
rect 78316 4274 78372 4284
rect 78876 4340 78932 4350
rect 78876 4246 78932 4284
rect 78764 4228 78820 4238
rect 78204 3666 78260 3678
rect 78204 3614 78206 3666
rect 78258 3614 78260 3666
rect 77532 3556 77588 3566
rect 77308 3554 77588 3556
rect 77308 3502 77534 3554
rect 77586 3502 77588 3554
rect 77308 3500 77588 3502
rect 77532 3490 77588 3500
rect 75740 3378 75796 3388
rect 75404 3332 75460 3342
rect 75404 800 75460 3276
rect 76300 3332 76356 3342
rect 76300 3238 76356 3276
rect 77420 812 77588 868
rect 77420 800 77476 812
rect 62440 200 62664 728
rect 63112 200 63336 728
rect 64456 200 64680 728
rect 64764 700 65492 756
rect 65800 200 66024 800
rect 67144 200 67368 800
rect 67816 200 68040 800
rect 69132 728 69384 800
rect 69160 200 69384 728
rect 70504 200 70728 800
rect 71176 200 71400 800
rect 72520 728 72772 800
rect 73864 728 74116 800
rect 75208 728 75460 800
rect 72520 200 72744 728
rect 73864 200 74088 728
rect 75208 200 75432 728
rect 75880 200 76104 800
rect 77224 728 77476 800
rect 77532 756 77588 812
rect 78204 756 78260 3614
rect 78764 800 78820 4172
rect 79548 4228 79604 4238
rect 79548 4134 79604 4172
rect 80556 3556 80612 4510
rect 81676 4564 81732 4844
rect 81676 4470 81732 4508
rect 83468 4564 83524 4574
rect 83468 4338 83524 4508
rect 83468 4286 83470 4338
rect 83522 4286 83524 4338
rect 83468 4274 83524 4286
rect 82348 4228 82404 4238
rect 82124 4226 82404 4228
rect 82124 4174 82350 4226
rect 82402 4174 82404 4226
rect 82124 4172 82404 4174
rect 81676 3666 81732 3678
rect 81676 3614 81678 3666
rect 81730 3614 81732 3666
rect 80892 3556 80948 3566
rect 80556 3554 80948 3556
rect 80556 3502 80894 3554
rect 80946 3502 80948 3554
rect 80556 3500 80948 3502
rect 80892 3490 80948 3500
rect 80220 3332 80276 3342
rect 80108 3330 80276 3332
rect 80108 3278 80222 3330
rect 80274 3278 80276 3330
rect 80108 3276 80276 3278
rect 80108 800 80164 3276
rect 80220 3266 80276 3276
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 81676 868 81732 3614
rect 80780 812 80948 868
rect 80780 800 80836 812
rect 77224 200 77448 728
rect 77532 700 78260 756
rect 78568 728 78820 800
rect 79912 728 80164 800
rect 80584 728 80836 800
rect 80892 756 80948 812
rect 81564 812 81732 868
rect 81564 756 81620 812
rect 82124 800 82180 4172
rect 82348 4162 82404 4172
rect 84140 3666 84196 27692
rect 84812 17668 84868 54348
rect 88508 54402 88564 54460
rect 89628 54516 89684 54526
rect 89628 54422 89684 54460
rect 88508 54350 88510 54402
rect 88562 54350 88564 54402
rect 86492 47460 86548 47470
rect 86492 24500 86548 47404
rect 87276 43538 87332 43550
rect 87276 43486 87278 43538
rect 87330 43486 87332 43538
rect 87276 43428 87332 43486
rect 87276 43362 87332 43372
rect 87836 43428 87892 43438
rect 87836 43334 87892 43372
rect 86492 24434 86548 24444
rect 86940 24948 86996 24958
rect 84812 17602 84868 17612
rect 86604 4452 86660 4462
rect 86492 4228 86548 4238
rect 86604 4228 86660 4396
rect 86492 4226 86660 4228
rect 86492 4174 86494 4226
rect 86546 4174 86660 4226
rect 86492 4172 86660 4174
rect 86492 4162 86548 4172
rect 84140 3614 84142 3666
rect 84194 3614 84196 3666
rect 84140 3602 84196 3614
rect 83468 3444 83524 3454
rect 83468 800 83524 3388
rect 85148 3444 85204 3454
rect 85148 3350 85204 3388
rect 86604 800 86660 4172
rect 86940 4226 86996 24892
rect 87948 4452 88004 4462
rect 87948 4358 88004 4396
rect 86940 4174 86942 4226
rect 86994 4174 86996 4226
rect 86940 4162 86996 4174
rect 88508 3666 88564 54350
rect 91532 51380 91588 64652
rect 93212 55860 93268 109228
rect 96636 109004 96900 109014
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96636 108938 96900 108948
rect 96636 107436 96900 107446
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96636 107370 96900 107380
rect 96636 105868 96900 105878
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96636 105802 96900 105812
rect 99820 105252 99876 116510
rect 100828 116340 100884 116350
rect 100828 116246 100884 116284
rect 100492 115554 100548 115566
rect 100492 115502 100494 115554
rect 100546 115502 100548 115554
rect 100492 115444 100548 115502
rect 100940 115556 100996 119200
rect 101612 116564 101668 116574
rect 100940 115490 100996 115500
rect 101052 115666 101108 115678
rect 101052 115614 101054 115666
rect 101106 115614 101108 115666
rect 100492 115378 100548 115388
rect 101052 115444 101108 115614
rect 101052 115378 101108 115388
rect 99820 105186 99876 105196
rect 100044 104580 100100 104590
rect 96636 104300 96900 104310
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96636 104234 96900 104244
rect 96636 102732 96900 102742
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96636 102666 96900 102676
rect 96636 101164 96900 101174
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96636 101098 96900 101108
rect 96636 99596 96900 99606
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96636 99530 96900 99540
rect 96636 98028 96900 98038
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96636 97962 96900 97972
rect 96636 96460 96900 96470
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96636 96394 96900 96404
rect 96636 94892 96900 94902
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96636 94826 96900 94836
rect 96636 93324 96900 93334
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96636 93258 96900 93268
rect 98252 92932 98308 92942
rect 96636 91756 96900 91766
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96636 91690 96900 91700
rect 96636 90188 96900 90198
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96636 90122 96900 90132
rect 96636 88620 96900 88630
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96636 88554 96900 88564
rect 96636 87052 96900 87062
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96636 86986 96900 86996
rect 96636 85484 96900 85494
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96636 85418 96900 85428
rect 96636 83916 96900 83926
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96636 83850 96900 83860
rect 96636 82348 96900 82358
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96636 82282 96900 82292
rect 96636 80780 96900 80790
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96636 80714 96900 80724
rect 96636 79212 96900 79222
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96636 79146 96900 79156
rect 96636 77644 96900 77654
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96636 77578 96900 77588
rect 96636 76076 96900 76086
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96636 76010 96900 76020
rect 96636 74508 96900 74518
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96636 74442 96900 74452
rect 96636 72940 96900 72950
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96636 72874 96900 72884
rect 96636 71372 96900 71382
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96636 71306 96900 71316
rect 96636 69804 96900 69814
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96636 69738 96900 69748
rect 96636 68236 96900 68246
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96636 68170 96900 68180
rect 96636 66668 96900 66678
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96636 66602 96900 66612
rect 96636 65100 96900 65110
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96636 65034 96900 65044
rect 96636 63532 96900 63542
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96636 63466 96900 63476
rect 98252 62356 98308 92876
rect 98252 62290 98308 62300
rect 96636 61964 96900 61974
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96636 61898 96900 61908
rect 98252 61796 98308 61806
rect 96636 60396 96900 60406
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96636 60330 96900 60340
rect 96636 58828 96900 58838
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96636 58762 96900 58772
rect 96636 57260 96900 57270
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96636 57194 96900 57204
rect 93212 55794 93268 55804
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 91532 51314 91588 51324
rect 92988 54740 93044 54750
rect 90188 50484 90244 50494
rect 90076 20580 90132 20590
rect 90076 20486 90132 20524
rect 90188 4340 90244 50428
rect 91532 47572 91588 47582
rect 91532 41972 91588 47516
rect 91532 41906 91588 41916
rect 91868 40964 91924 40974
rect 91756 22260 91812 22270
rect 91196 22258 91812 22260
rect 91196 22206 91758 22258
rect 91810 22206 91812 22258
rect 91196 22204 91812 22206
rect 90636 21476 90692 21486
rect 90636 21382 90692 21420
rect 91196 21026 91252 22204
rect 91756 22194 91812 22204
rect 91308 21588 91364 21598
rect 91308 21494 91364 21532
rect 91196 20974 91198 21026
rect 91250 20974 91252 21026
rect 91196 20962 91252 20974
rect 90524 20804 90580 20814
rect 90524 20578 90580 20748
rect 91532 20804 91588 20814
rect 91532 20710 91588 20748
rect 90524 20526 90526 20578
rect 90578 20526 90580 20578
rect 90524 4564 90580 20526
rect 91868 20188 91924 40908
rect 92092 22146 92148 22158
rect 92092 22094 92094 22146
rect 92146 22094 92148 22146
rect 91980 21700 92036 21710
rect 92092 21700 92148 22094
rect 91980 21698 92148 21700
rect 91980 21646 91982 21698
rect 92034 21646 92148 21698
rect 91980 21644 92148 21646
rect 91980 21634 92036 21644
rect 92204 20804 92260 20814
rect 92204 20580 92260 20748
rect 92316 20692 92372 20702
rect 92316 20598 92372 20636
rect 92204 20514 92260 20524
rect 91868 20132 92036 20188
rect 90524 4498 90580 4508
rect 90188 4274 90244 4284
rect 88508 3614 88510 3666
rect 88562 3614 88564 3666
rect 88508 3556 88564 3614
rect 91980 3666 92036 20132
rect 92652 4452 92708 4462
rect 92540 4228 92596 4238
rect 92652 4228 92708 4396
rect 92540 4226 92708 4228
rect 92540 4174 92542 4226
rect 92594 4174 92708 4226
rect 92540 4172 92708 4174
rect 92540 4162 92596 4172
rect 91980 3614 91982 3666
rect 92034 3614 92036 3666
rect 91980 3602 92036 3614
rect 88508 3490 88564 3500
rect 89964 3556 90020 3566
rect 89964 3462 90020 3500
rect 89068 3444 89124 3454
rect 88844 3442 89124 3444
rect 88844 3390 89070 3442
rect 89122 3390 89124 3442
rect 88844 3388 89124 3390
rect 88844 800 88900 3388
rect 89068 3378 89124 3388
rect 91308 3444 91364 3454
rect 91308 800 91364 3388
rect 92652 800 92708 4172
rect 92988 4226 93044 54684
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 96636 47852 96900 47862
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 96636 46284 96900 46294
rect 94892 46228 94948 46238
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 94892 33572 94948 46172
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 95676 35700 95732 35710
rect 95676 34692 95732 35644
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 95676 34626 95732 34636
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 94892 33506 94948 33516
rect 95228 32452 95284 32462
rect 93100 21476 93156 21486
rect 93100 20914 93156 21420
rect 94108 21476 94164 21486
rect 94108 21382 94164 21420
rect 95004 21476 95060 21486
rect 93100 20862 93102 20914
rect 93154 20862 93156 20914
rect 93100 20692 93156 20862
rect 93100 20626 93156 20636
rect 93996 4452 94052 4462
rect 93996 4358 94052 4396
rect 95004 4340 95060 21420
rect 95228 20804 95284 32396
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 95228 20738 95284 20748
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 98252 6804 98308 61740
rect 100044 52052 100100 104524
rect 101612 54292 101668 116508
rect 106876 116562 106932 119200
rect 106876 116510 106878 116562
rect 106930 116510 106932 116562
rect 106876 116340 106932 116510
rect 106876 116274 106932 116284
rect 107660 116562 107716 116574
rect 107660 116510 107662 116562
rect 107714 116510 107716 116562
rect 101724 115556 101780 115566
rect 101724 115462 101780 115500
rect 103292 115556 103348 115566
rect 103292 62580 103348 115500
rect 106652 107716 106708 107726
rect 103292 62514 103348 62524
rect 104972 74228 105028 74238
rect 103516 55524 103572 55534
rect 101612 54226 101668 54236
rect 101836 55300 101892 55310
rect 100044 51986 100100 51996
rect 100268 51156 100324 51166
rect 100268 14308 100324 51100
rect 100828 43428 100884 43438
rect 100828 41188 100884 43372
rect 101836 43428 101892 55244
rect 101836 43362 101892 43372
rect 100828 41122 100884 41132
rect 100268 14242 100324 14252
rect 101836 40404 101892 40414
rect 101836 12068 101892 40348
rect 101836 12002 101892 12012
rect 103292 37828 103348 37838
rect 98252 6738 98308 6748
rect 100268 9268 100324 9278
rect 92988 4174 92990 4226
rect 93042 4174 93044 4226
rect 92988 4162 93044 4174
rect 94780 4338 95060 4340
rect 94780 4286 95006 4338
rect 95058 4286 95060 4338
rect 94780 4284 95060 4286
rect 94780 3666 94836 4284
rect 95004 4274 95060 4284
rect 96348 5908 96404 5918
rect 94780 3614 94782 3666
rect 94834 3614 94836 3666
rect 94780 3602 94836 3614
rect 95676 4226 95732 4238
rect 95676 4174 95678 4226
rect 95730 4174 95732 4226
rect 92988 3444 93044 3454
rect 92988 3350 93044 3388
rect 94892 812 95060 868
rect 94892 800 94948 812
rect 78568 200 78792 728
rect 79912 200 80136 728
rect 80584 200 80808 728
rect 80892 700 81620 756
rect 81928 728 82180 800
rect 83272 728 83524 800
rect 81928 200 82152 728
rect 83272 200 83496 728
rect 83944 200 84168 800
rect 85288 200 85512 800
rect 86604 728 86856 800
rect 86632 200 86856 728
rect 87976 200 88200 800
rect 88648 728 88900 800
rect 88648 200 88872 728
rect 89992 200 90216 800
rect 91308 728 91560 800
rect 92652 728 92904 800
rect 91336 200 91560 728
rect 92680 200 92904 728
rect 93352 200 93576 800
rect 94696 728 94948 800
rect 95004 756 95060 812
rect 95676 756 95732 4174
rect 96348 3666 96404 5852
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 99148 5012 99204 5022
rect 99148 4918 99204 4956
rect 99932 5012 99988 5022
rect 99484 4898 99540 4910
rect 99484 4846 99486 4898
rect 99538 4846 99540 4898
rect 98028 4452 98084 4462
rect 97916 4228 97972 4238
rect 98028 4228 98084 4396
rect 99372 4452 99428 4462
rect 99372 4358 99428 4396
rect 97916 4226 98084 4228
rect 97916 4174 97918 4226
rect 97970 4174 98084 4226
rect 97916 4172 98084 4174
rect 97916 4162 97972 4172
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 96348 3614 96350 3666
rect 96402 3614 96404 3666
rect 96348 3602 96404 3614
rect 95900 3444 95956 3454
rect 96012 3444 96068 3454
rect 95900 3442 96012 3444
rect 95900 3390 95902 3442
rect 95954 3390 96012 3442
rect 95900 3388 96012 3390
rect 95900 3378 95956 3388
rect 94696 200 94920 728
rect 95004 700 95732 756
rect 96012 800 96068 3388
rect 97356 3444 97412 3454
rect 97356 3350 97412 3388
rect 98028 800 98084 4172
rect 98364 4340 98420 4350
rect 98364 4226 98420 4284
rect 98364 4174 98366 4226
rect 98418 4174 98420 4226
rect 98364 4162 98420 4174
rect 99484 3556 99540 4846
rect 99932 4898 99988 4956
rect 99932 4846 99934 4898
rect 99986 4846 99988 4898
rect 99932 4340 99988 4846
rect 99932 4274 99988 4284
rect 100268 4226 100324 9212
rect 101388 4898 101444 4910
rect 101388 4846 101390 4898
rect 101442 4846 101444 4898
rect 101388 4564 101444 4846
rect 101388 4498 101444 4508
rect 103292 4564 103348 37772
rect 103516 37828 103572 55468
rect 104972 55188 105028 74172
rect 106652 60228 106708 107660
rect 107660 64708 107716 116510
rect 108668 116340 108724 116350
rect 108668 116246 108724 116284
rect 108668 115892 108724 115902
rect 108780 115892 108836 119200
rect 108668 115890 108836 115892
rect 108668 115838 108670 115890
rect 108722 115838 108836 115890
rect 108668 115836 108836 115838
rect 108668 115826 108724 115836
rect 108780 115780 108836 115836
rect 108780 115714 108836 115724
rect 110124 115780 110180 115790
rect 110124 115686 110180 115724
rect 110348 115780 110404 119200
rect 110908 119308 111412 119364
rect 111496 119336 111720 119800
rect 110908 116562 110964 119308
rect 111356 119140 111412 119308
rect 111468 119200 111720 119336
rect 112168 119200 112392 119800
rect 113512 119200 113736 119800
rect 114856 119336 115080 119800
rect 114828 119200 115080 119336
rect 115528 119200 115752 119800
rect 116872 119336 117096 119800
rect 116844 119200 117096 119336
rect 118216 119200 118440 119800
rect 119560 119200 119784 119800
rect 111468 119140 111524 119200
rect 111356 119084 111524 119140
rect 110908 116510 110910 116562
rect 110962 116510 110964 116562
rect 110908 116340 110964 116510
rect 111804 116564 111860 116574
rect 111804 116470 111860 116508
rect 114828 116562 114884 119200
rect 114828 116510 114830 116562
rect 114882 116510 114884 116562
rect 110908 116274 110964 116284
rect 112812 116340 112868 116350
rect 112812 116246 112868 116284
rect 114828 116340 114884 116510
rect 115724 116564 115780 116574
rect 115724 116470 115780 116508
rect 114828 116274 114884 116284
rect 116508 116340 116564 116350
rect 116508 116246 116564 116284
rect 111996 116060 112260 116070
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 111996 115994 112260 116004
rect 110348 115714 110404 115724
rect 111244 115780 111300 115790
rect 111244 115686 111300 115724
rect 112364 115668 112420 115678
rect 116172 115668 116228 115678
rect 112364 115666 112644 115668
rect 112364 115614 112366 115666
rect 112418 115614 112644 115666
rect 112364 115612 112644 115614
rect 112364 115602 112420 115612
rect 109116 115556 109172 115566
rect 109116 115462 109172 115500
rect 110796 114884 110852 114894
rect 110796 114790 110852 114828
rect 112588 114884 112644 115612
rect 116172 115666 116676 115668
rect 116172 115614 116174 115666
rect 116226 115614 116676 115666
rect 116172 115612 116676 115614
rect 116172 115602 116228 115612
rect 115500 115556 115556 115566
rect 115500 115462 115556 115500
rect 115836 115332 115892 115342
rect 115500 115220 115556 115230
rect 111996 114492 112260 114502
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 111996 114426 112260 114436
rect 111996 112924 112260 112934
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 111996 112858 112260 112868
rect 111996 111356 112260 111366
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 111996 111290 112260 111300
rect 111996 109788 112260 109798
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 111996 109722 112260 109732
rect 111996 108220 112260 108230
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 111996 108154 112260 108164
rect 111996 106652 112260 106662
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 111996 106586 112260 106596
rect 111996 105084 112260 105094
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 111996 105018 112260 105028
rect 111996 103516 112260 103526
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 111996 103450 112260 103460
rect 111996 101948 112260 101958
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 111996 101882 112260 101892
rect 111996 100380 112260 100390
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 111996 100314 112260 100324
rect 111996 98812 112260 98822
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 111996 98746 112260 98756
rect 111996 97244 112260 97254
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 111996 97178 112260 97188
rect 111996 95676 112260 95686
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 111996 95610 112260 95620
rect 111996 94108 112260 94118
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 111996 94042 112260 94052
rect 111996 92540 112260 92550
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 111996 92474 112260 92484
rect 111996 90972 112260 90982
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 111996 90906 112260 90916
rect 111996 89404 112260 89414
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 111996 89338 112260 89348
rect 111996 87836 112260 87846
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 111996 87770 112260 87780
rect 111996 86268 112260 86278
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 111996 86202 112260 86212
rect 111996 84700 112260 84710
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 111996 84634 112260 84644
rect 111996 83132 112260 83142
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 111996 83066 112260 83076
rect 111996 81564 112260 81574
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 111996 81498 112260 81508
rect 111996 79996 112260 80006
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 111996 79930 112260 79940
rect 111996 78428 112260 78438
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 111996 78362 112260 78372
rect 111996 76860 112260 76870
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 111996 76794 112260 76804
rect 111996 75292 112260 75302
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 111996 75226 112260 75236
rect 111996 73724 112260 73734
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 111996 73658 112260 73668
rect 111996 72156 112260 72166
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 111996 72090 112260 72100
rect 111996 70588 112260 70598
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 111996 70522 112260 70532
rect 111996 69020 112260 69030
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 111996 68954 112260 68964
rect 111996 67452 112260 67462
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 111996 67386 112260 67396
rect 111996 65884 112260 65894
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 111996 65818 112260 65828
rect 107660 64642 107716 64652
rect 108332 64820 108388 64830
rect 108332 63252 108388 64764
rect 111996 64316 112260 64326
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 111996 64250 112260 64260
rect 108332 63186 108388 63196
rect 111996 62748 112260 62758
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 111996 62682 112260 62692
rect 111996 61180 112260 61190
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 111996 61114 112260 61124
rect 106652 60162 106708 60172
rect 111996 59612 112260 59622
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 111996 59546 112260 59556
rect 108332 59332 108388 59342
rect 108332 58548 108388 59276
rect 108332 58482 108388 58492
rect 104972 55122 105028 55132
rect 110236 58324 110292 58334
rect 103516 37762 103572 37772
rect 104972 53508 105028 53518
rect 104972 5796 105028 53452
rect 108220 52836 108276 52846
rect 108220 46564 108276 52780
rect 108220 46498 108276 46508
rect 108332 47236 108388 47246
rect 104972 5730 105028 5740
rect 103292 4498 103348 4508
rect 104300 5012 104356 5022
rect 104300 4562 104356 4956
rect 104300 4510 104302 4562
rect 104354 4510 104356 4562
rect 101164 4450 101220 4462
rect 101164 4398 101166 4450
rect 101218 4398 101220 4450
rect 100940 4340 100996 4350
rect 101164 4340 101220 4398
rect 103516 4452 103572 4462
rect 103516 4358 103572 4396
rect 103852 4450 103908 4462
rect 103852 4398 103854 4450
rect 103906 4398 103908 4450
rect 101724 4340 101780 4350
rect 101164 4338 101780 4340
rect 101164 4286 101726 4338
rect 101778 4286 101780 4338
rect 101164 4284 101780 4286
rect 100940 4246 100996 4284
rect 101724 4274 101780 4284
rect 100268 4174 100270 4226
rect 100322 4174 100324 4226
rect 99820 3556 99876 3566
rect 99484 3554 99876 3556
rect 99484 3502 99822 3554
rect 99874 3502 99876 3554
rect 99484 3500 99876 3502
rect 99820 3490 99876 3500
rect 100268 3556 100324 4174
rect 102396 4226 102452 4238
rect 102396 4174 102398 4226
rect 102450 4174 102452 4226
rect 100492 3668 100548 3678
rect 100268 3490 100324 3500
rect 100380 3666 100548 3668
rect 100380 3614 100494 3666
rect 100546 3614 100548 3666
rect 100380 3612 100548 3614
rect 99596 812 99764 868
rect 99596 800 99652 812
rect 96012 728 96264 800
rect 96040 200 96264 728
rect 96712 200 96936 800
rect 98028 728 98280 800
rect 98056 200 98280 728
rect 99400 728 99652 800
rect 99708 756 99764 812
rect 100380 756 100436 3612
rect 100492 3602 100548 3612
rect 100940 3444 100996 3454
rect 100940 800 100996 3388
rect 101724 3444 101780 3454
rect 101724 3350 101780 3388
rect 101612 812 101780 868
rect 101612 800 101668 812
rect 99400 200 99624 728
rect 99708 700 100436 756
rect 100744 728 100996 800
rect 101416 728 101668 800
rect 101724 756 101780 812
rect 102396 756 102452 4174
rect 102956 3668 103012 3678
rect 102620 3556 102676 3566
rect 102620 3462 102676 3500
rect 102956 800 103012 3612
rect 103852 3554 103908 4398
rect 104300 4452 104356 4510
rect 104300 4386 104356 4396
rect 104412 3668 104468 3678
rect 104412 3574 104468 3612
rect 108332 3668 108388 47180
rect 110236 35252 110292 58268
rect 111996 58044 112260 58054
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 111996 57978 112260 57988
rect 111996 56476 112260 56486
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 111996 56410 112260 56420
rect 111996 54908 112260 54918
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 111996 54842 112260 54852
rect 111996 53340 112260 53350
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 111996 53274 112260 53284
rect 111996 51772 112260 51782
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 111996 51706 112260 51716
rect 111996 50204 112260 50214
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 111996 50138 112260 50148
rect 111996 48636 112260 48646
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 111996 48570 112260 48580
rect 111996 47068 112260 47078
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 111996 47002 112260 47012
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 110236 35186 110292 35196
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 110012 34020 110068 34030
rect 110012 21588 110068 33964
rect 112588 33572 112644 114828
rect 114380 114884 114436 114894
rect 114380 114790 114436 114828
rect 115164 114884 115220 114894
rect 115164 114790 115220 114828
rect 115500 113986 115556 115164
rect 115836 114994 115892 115276
rect 116620 115108 116676 115612
rect 116844 115332 116900 119200
rect 117852 118244 117908 118254
rect 117516 116226 117572 116238
rect 117516 116174 117518 116226
rect 117570 116174 117572 116226
rect 116956 115668 117012 115678
rect 117516 115668 117572 116174
rect 117852 115778 117908 118188
rect 117852 115726 117854 115778
rect 117906 115726 117908 115778
rect 117852 115714 117908 115726
rect 118188 116564 118244 116574
rect 116956 115666 117572 115668
rect 116956 115614 116958 115666
rect 117010 115614 117572 115666
rect 116956 115612 117572 115614
rect 116956 115602 117012 115612
rect 116844 115266 116900 115276
rect 116620 115052 117124 115108
rect 115836 114942 115838 114994
rect 115890 114942 115892 114994
rect 115836 114930 115892 114942
rect 116284 114996 116340 115006
rect 116284 114324 116340 114940
rect 117068 114770 117124 115052
rect 117068 114718 117070 114770
rect 117122 114718 117124 114770
rect 117068 114706 117124 114718
rect 117180 114548 117236 115612
rect 116284 114258 116340 114268
rect 116396 114492 117236 114548
rect 117292 114882 117348 114894
rect 117292 114830 117294 114882
rect 117346 114830 117348 114882
rect 115500 113934 115502 113986
rect 115554 113934 115556 113986
rect 115500 113922 115556 113934
rect 116172 114098 116228 114110
rect 116172 114046 116174 114098
rect 116226 114046 116228 114098
rect 116172 113986 116228 114046
rect 116172 113934 116174 113986
rect 116226 113934 116228 113986
rect 116172 113922 116228 113934
rect 115164 110964 115220 110974
rect 115500 110964 115556 110974
rect 115164 110962 115500 110964
rect 115164 110910 115166 110962
rect 115218 110910 115500 110962
rect 115164 110908 115500 110910
rect 115164 110898 115220 110908
rect 114940 109284 114996 109294
rect 114940 109190 114996 109228
rect 114940 107716 114996 107726
rect 114940 107622 114996 107660
rect 114492 106260 114548 106270
rect 114492 106166 114548 106204
rect 114940 106260 114996 106270
rect 114940 106166 114996 106204
rect 114940 104580 114996 104590
rect 114940 104486 114996 104524
rect 114828 102452 114884 102462
rect 114828 102358 114884 102396
rect 114492 99988 114548 99998
rect 114940 99988 114996 99998
rect 114492 99986 114996 99988
rect 114492 99934 114494 99986
rect 114546 99934 114942 99986
rect 114994 99934 114996 99986
rect 114492 99932 114996 99934
rect 114492 99876 114548 99932
rect 114940 99922 114996 99932
rect 114492 99810 114548 99820
rect 114940 95282 114996 95294
rect 114940 95230 114942 95282
rect 114994 95230 114996 95282
rect 114492 95172 114548 95182
rect 114940 95172 114996 95230
rect 114492 95170 114996 95172
rect 114492 95118 114494 95170
rect 114546 95118 114996 95170
rect 114492 95116 114996 95118
rect 114492 94276 114548 95116
rect 114828 94612 114884 94622
rect 114828 94518 114884 94556
rect 114492 94210 114548 94220
rect 114380 92932 114436 92942
rect 114380 92838 114436 92876
rect 114940 92932 114996 92942
rect 114940 92838 114996 92876
rect 115388 89906 115444 89918
rect 115388 89854 115390 89906
rect 115442 89854 115444 89906
rect 115388 89572 115444 89854
rect 115388 89506 115444 89516
rect 114940 87332 114996 87342
rect 114940 87238 114996 87276
rect 114380 86660 114436 86670
rect 114380 86566 114436 86604
rect 114940 86660 114996 86670
rect 114940 86566 114996 86604
rect 114492 85092 114548 85102
rect 114940 85092 114996 85102
rect 114492 85090 114996 85092
rect 114492 85038 114494 85090
rect 114546 85038 114942 85090
rect 114994 85038 114996 85090
rect 114492 85036 114996 85038
rect 114492 84868 114548 85036
rect 114940 85026 114996 85036
rect 114492 84802 114548 84812
rect 115388 83634 115444 83646
rect 115388 83582 115390 83634
rect 115442 83582 115444 83634
rect 115388 83524 115444 83582
rect 115388 83458 115444 83468
rect 114828 79380 114884 79390
rect 114828 79286 114884 79324
rect 114828 77812 114884 77822
rect 114828 77718 114884 77756
rect 114380 75684 114436 75694
rect 114380 75590 114436 75628
rect 114940 75684 114996 75694
rect 114940 75590 114996 75628
rect 114828 74228 114884 74238
rect 114828 74134 114884 74172
rect 115500 70418 115556 110908
rect 115836 110850 115892 110862
rect 115836 110798 115838 110850
rect 115890 110798 115892 110850
rect 115836 110404 115892 110798
rect 115836 110338 115892 110348
rect 116284 109506 116340 109518
rect 116284 109454 116286 109506
rect 116338 109454 116340 109506
rect 116284 109284 116340 109454
rect 116284 109218 116340 109228
rect 116284 107938 116340 107950
rect 116284 107886 116286 107938
rect 116338 107886 116340 107938
rect 116284 107716 116340 107886
rect 116284 107650 116340 107660
rect 115836 106146 115892 106158
rect 115836 106094 115838 106146
rect 115890 106094 115892 106146
rect 115836 105700 115892 106094
rect 115836 105634 115892 105644
rect 116284 104802 116340 104814
rect 116284 104750 116286 104802
rect 116338 104750 116340 104802
rect 116284 104356 116340 104750
rect 116284 104290 116340 104300
rect 116396 102508 116452 114492
rect 116620 114324 116676 114334
rect 116620 111076 116676 114268
rect 117068 114324 117124 114362
rect 117292 114324 117348 114830
rect 117124 114268 117348 114324
rect 117740 114884 117796 114894
rect 117068 114258 117124 114268
rect 116732 113988 116788 113998
rect 116732 113986 117012 113988
rect 116732 113934 116734 113986
rect 116786 113934 117012 113986
rect 116732 113932 117012 113934
rect 116732 113874 116788 113932
rect 116732 113822 116734 113874
rect 116786 113822 116788 113874
rect 116732 113810 116788 113822
rect 116620 111020 116788 111076
rect 116508 110964 116564 110974
rect 116564 110908 116676 110964
rect 116508 110898 116564 110908
rect 116620 110850 116676 110908
rect 116620 110798 116622 110850
rect 116674 110798 116676 110850
rect 116620 110786 116676 110798
rect 116172 102452 116452 102508
rect 116060 102226 116116 102238
rect 116060 102174 116062 102226
rect 116114 102174 116116 102226
rect 116060 102116 116116 102174
rect 116060 102050 116116 102060
rect 115836 99874 115892 99886
rect 115836 99822 115838 99874
rect 115890 99822 115892 99874
rect 115836 99652 115892 99822
rect 115836 99586 115892 99596
rect 115836 95170 115892 95182
rect 115836 95118 115838 95170
rect 115890 95118 115892 95170
rect 115836 94948 115892 95118
rect 115836 94882 115892 94892
rect 116060 94386 116116 94398
rect 116060 94334 116062 94386
rect 116114 94334 116116 94386
rect 116060 94276 116116 94334
rect 116060 94210 116116 94220
rect 115836 93042 115892 93054
rect 115836 92990 115838 93042
rect 115890 92990 115892 93042
rect 115836 92932 115892 92990
rect 115836 92866 115892 92876
rect 116172 90748 116228 102452
rect 116060 90692 116228 90748
rect 115948 89794 116004 89806
rect 115948 89742 115950 89794
rect 116002 89742 116004 89794
rect 115948 89684 116004 89742
rect 115836 86770 115892 86782
rect 115836 86718 115838 86770
rect 115890 86718 115892 86770
rect 115836 86212 115892 86718
rect 115836 86146 115892 86156
rect 115836 85202 115892 85214
rect 115836 85150 115838 85202
rect 115890 85150 115892 85202
rect 115836 84868 115892 85150
rect 115836 84802 115892 84812
rect 115948 73108 116004 89628
rect 116060 78988 116116 90692
rect 116284 87556 116340 87566
rect 116284 87462 116340 87500
rect 116732 83636 116788 111020
rect 116844 109284 116900 109294
rect 116844 109190 116900 109228
rect 116844 107716 116900 107726
rect 116844 107622 116900 107660
rect 116844 104578 116900 104590
rect 116844 104526 116846 104578
rect 116898 104526 116900 104578
rect 116844 104356 116900 104526
rect 116844 104290 116900 104300
rect 116956 102508 117012 113932
rect 116956 102452 117572 102508
rect 117068 102116 117124 102126
rect 117068 102022 117124 102060
rect 117068 94276 117124 94286
rect 117068 94182 117124 94220
rect 116956 89684 117012 89694
rect 116956 89590 117012 89628
rect 116844 87556 116900 87566
rect 116844 87442 116900 87500
rect 116844 87390 116846 87442
rect 116898 87390 116900 87442
rect 116844 86884 116900 87390
rect 116844 86818 116900 86828
rect 116732 83580 117348 83636
rect 116172 83522 116228 83534
rect 116172 83470 116174 83522
rect 116226 83470 116228 83522
rect 116172 83412 116228 83470
rect 116172 83346 116228 83356
rect 116732 82962 116788 83580
rect 117292 83522 117348 83580
rect 117292 83470 117294 83522
rect 117346 83470 117348 83522
rect 117292 83458 117348 83470
rect 117068 83412 117124 83422
rect 117068 83318 117124 83356
rect 116732 82910 116734 82962
rect 116786 82910 116788 82962
rect 116732 82898 116788 82910
rect 117292 79940 117348 79950
rect 117292 79714 117348 79884
rect 117292 79662 117294 79714
rect 117346 79662 117348 79714
rect 117292 79650 117348 79662
rect 117516 78988 117572 102452
rect 116060 78932 116564 78988
rect 116060 75570 116116 75582
rect 116060 75518 116062 75570
rect 116114 75518 116116 75570
rect 116060 75460 116116 75518
rect 116060 75394 116116 75404
rect 116172 74004 116228 74014
rect 116172 73910 116228 73948
rect 115948 73052 116452 73108
rect 116396 71092 116452 73052
rect 116060 71036 116452 71092
rect 115500 70366 115502 70418
rect 115554 70366 115556 70418
rect 114380 69412 114436 69422
rect 114380 69318 114436 69356
rect 114940 69412 114996 69422
rect 114940 69318 114996 69356
rect 115164 68852 115220 68862
rect 114492 68628 114548 68638
rect 114156 68626 114548 68628
rect 114156 68574 114494 68626
rect 114546 68574 114548 68626
rect 114156 68572 114548 68574
rect 114044 68516 114100 68526
rect 114156 68516 114212 68572
rect 114492 68562 114548 68572
rect 114044 68514 114212 68516
rect 114044 68462 114046 68514
rect 114098 68462 114212 68514
rect 114044 68460 114212 68462
rect 114044 68450 114100 68460
rect 114156 67284 114212 68460
rect 114156 67218 114212 67228
rect 113932 66948 113988 66958
rect 112700 66164 112756 66174
rect 112700 65604 112756 66108
rect 113484 66164 113540 66174
rect 113484 66070 113540 66108
rect 113932 65716 113988 66892
rect 114380 66946 114436 66958
rect 114380 66894 114382 66946
rect 114434 66894 114436 66946
rect 114380 66500 114436 66894
rect 115164 66946 115220 68796
rect 115500 68852 115556 70366
rect 115948 70420 116004 70430
rect 115500 68786 115556 68796
rect 115836 69522 115892 69534
rect 115836 69470 115838 69522
rect 115890 69470 115892 69522
rect 115836 68740 115892 69470
rect 115836 68674 115892 68684
rect 115612 68514 115668 68526
rect 115612 68462 115614 68514
rect 115666 68462 115668 68514
rect 115164 66894 115166 66946
rect 115218 66894 115220 66946
rect 115164 66882 115220 66894
rect 115500 67954 115556 67966
rect 115500 67902 115502 67954
rect 115554 67902 115556 67954
rect 114380 66444 115220 66500
rect 114156 66276 114212 66286
rect 114156 66182 114212 66220
rect 115052 66276 115108 66286
rect 115164 66276 115220 66444
rect 115388 66276 115444 66286
rect 115164 66274 115444 66276
rect 115164 66222 115390 66274
rect 115442 66222 115444 66274
rect 115164 66220 115444 66222
rect 115052 66182 115108 66220
rect 114380 66052 114436 66062
rect 114380 66050 114996 66052
rect 114380 65998 114382 66050
rect 114434 65998 114996 66050
rect 114380 65996 114996 65998
rect 114380 65986 114436 65996
rect 113932 65584 113988 65660
rect 114492 65716 114548 65726
rect 114940 65716 114996 65996
rect 114940 65660 115332 65716
rect 112700 65538 112756 65548
rect 114492 65490 114548 65660
rect 115276 65602 115332 65660
rect 115276 65550 115278 65602
rect 115330 65550 115332 65602
rect 115276 65538 115332 65550
rect 114492 65438 114494 65490
rect 114546 65438 114548 65490
rect 114492 65426 114548 65438
rect 114828 64820 114884 64830
rect 114828 64726 114884 64764
rect 114828 63364 114884 63374
rect 114828 63250 114884 63308
rect 114828 63198 114830 63250
rect 114882 63198 114884 63250
rect 114828 63186 114884 63198
rect 114828 62132 114884 62142
rect 114828 61682 114884 62076
rect 114828 61630 114830 61682
rect 114882 61630 114884 61682
rect 114828 61618 114884 61630
rect 114940 60674 114996 60686
rect 114940 60622 114942 60674
rect 114994 60622 114996 60674
rect 114940 60004 114996 60622
rect 114940 59938 114996 59948
rect 114940 59778 114996 59790
rect 114940 59726 114942 59778
rect 114994 59726 114996 59778
rect 114940 59444 114996 59726
rect 115276 59780 115332 59790
rect 115276 59686 115332 59724
rect 114940 59378 114996 59388
rect 114828 58548 114884 58558
rect 114828 58454 114884 58492
rect 114492 56196 114548 56206
rect 114492 56102 114548 56140
rect 114940 56196 114996 56206
rect 114940 56082 114996 56140
rect 114940 56030 114942 56082
rect 114994 56030 114996 56082
rect 114940 56018 114996 56030
rect 114380 55300 114436 55310
rect 114380 55074 114436 55244
rect 114940 55300 114996 55310
rect 114940 55206 114996 55244
rect 114380 55022 114382 55074
rect 114434 55022 114436 55074
rect 114380 54628 114436 55022
rect 114380 54562 114436 54572
rect 114940 52836 114996 52846
rect 114940 52742 114996 52780
rect 115388 45332 115444 66220
rect 115500 66052 115556 67902
rect 115612 67396 115668 68462
rect 115612 67330 115668 67340
rect 115948 67172 116004 70364
rect 115612 66836 115668 66846
rect 115612 66164 115668 66780
rect 115612 66070 115668 66108
rect 115500 65986 115556 65996
rect 115948 65940 116004 67116
rect 116060 66164 116116 71036
rect 116508 70420 116564 78932
rect 117292 78932 117572 78988
rect 117180 78596 117236 78606
rect 117180 78146 117236 78540
rect 117180 78094 117182 78146
rect 117234 78094 117236 78146
rect 117180 78082 117236 78094
rect 117068 74004 117124 74014
rect 117068 73444 117124 73948
rect 117068 73378 117124 73388
rect 116508 70354 116564 70364
rect 117068 69186 117124 69198
rect 117068 69134 117070 69186
rect 117122 69134 117124 69186
rect 116396 68852 116452 68862
rect 116396 68738 116452 68796
rect 116396 68686 116398 68738
rect 116450 68686 116452 68738
rect 116396 68674 116452 68686
rect 116956 68740 117012 68750
rect 117068 68740 117124 69134
rect 116956 68738 117124 68740
rect 116956 68686 116958 68738
rect 117010 68686 117124 68738
rect 116956 68684 117124 68686
rect 116172 67842 116228 67854
rect 116172 67790 116174 67842
rect 116226 67790 116228 67842
rect 116172 67228 116228 67790
rect 116172 67172 116900 67228
rect 116844 66612 116900 67172
rect 116956 66836 117012 68684
rect 117180 68402 117236 68414
rect 117180 68350 117182 68402
rect 117234 68350 117236 68402
rect 117068 67618 117124 67630
rect 117068 67566 117070 67618
rect 117122 67566 117124 67618
rect 117068 67228 117124 67566
rect 117180 67508 117236 68350
rect 117292 67620 117348 78932
rect 117516 68402 117572 68414
rect 117516 68350 117518 68402
rect 117570 68350 117572 68402
rect 117404 67844 117460 67854
rect 117516 67844 117572 68350
rect 117404 67842 117572 67844
rect 117404 67790 117406 67842
rect 117458 67790 117572 67842
rect 117404 67788 117572 67790
rect 117404 67778 117460 67788
rect 117292 67564 117572 67620
rect 117180 67452 117460 67508
rect 117068 67172 117348 67228
rect 117292 67170 117348 67172
rect 117292 67118 117294 67170
rect 117346 67118 117348 67170
rect 117292 67106 117348 67118
rect 117404 67172 117460 67452
rect 116956 66770 117012 66780
rect 116844 66556 117124 66612
rect 116060 66032 116116 66108
rect 117068 66162 117124 66556
rect 117404 66276 117460 67116
rect 117068 66110 117070 66162
rect 117122 66110 117124 66162
rect 117068 66098 117124 66110
rect 117292 66164 117348 66174
rect 117404 66144 117460 66220
rect 117292 65940 117348 66108
rect 117292 65884 117460 65940
rect 115948 65874 116004 65884
rect 117404 65378 117460 65884
rect 117404 65326 117406 65378
rect 117458 65326 117460 65378
rect 117404 65314 117460 65326
rect 116172 65156 116228 65166
rect 116172 64594 116228 65100
rect 116956 65156 117012 65166
rect 116956 64818 117012 65100
rect 116956 64766 116958 64818
rect 117010 64766 117012 64818
rect 116956 64754 117012 64766
rect 116172 64542 116174 64594
rect 116226 64542 116228 64594
rect 116172 64530 116228 64542
rect 116172 63026 116228 63038
rect 116172 62974 116174 63026
rect 116226 62974 116228 63026
rect 116172 62692 116228 62974
rect 116172 62626 116228 62636
rect 117068 62914 117124 62926
rect 117068 62862 117070 62914
rect 117122 62862 117124 62914
rect 117068 62692 117124 62862
rect 117068 62626 117124 62636
rect 116172 61458 116228 61470
rect 116172 61406 116174 61458
rect 116226 61406 116228 61458
rect 116172 61348 116228 61406
rect 116172 61282 116228 61292
rect 117068 61348 117124 61358
rect 117068 61254 117124 61292
rect 116284 60898 116340 60910
rect 116284 60846 116286 60898
rect 116338 60846 116340 60898
rect 116284 60676 116340 60846
rect 116284 60610 116340 60620
rect 116844 60676 116900 60686
rect 116844 60582 116900 60620
rect 115836 59780 115892 59790
rect 115836 59332 115892 59724
rect 115836 59266 115892 59276
rect 116172 58322 116228 58334
rect 116172 58270 116174 58322
rect 116226 58270 116228 58322
rect 116172 57988 116228 58270
rect 116172 57922 116228 57932
rect 117068 58210 117124 58222
rect 117068 58158 117070 58210
rect 117122 58158 117124 58210
rect 117068 57988 117124 58158
rect 117516 57988 117572 67564
rect 117740 67228 117796 114828
rect 118076 112644 118132 112654
rect 118076 112550 118132 112588
rect 118076 111524 118132 111534
rect 118076 111430 118132 111468
rect 118076 106820 118132 106830
rect 118076 106726 118132 106764
rect 118076 101666 118132 101678
rect 118076 101614 118078 101666
rect 118130 101614 118132 101666
rect 118076 100996 118132 101614
rect 118076 100930 118132 100940
rect 118076 96962 118132 96974
rect 118076 96910 118078 96962
rect 118130 96910 118132 96962
rect 118076 96292 118132 96910
rect 118076 96226 118132 96236
rect 118076 82850 118132 82862
rect 118076 82798 118078 82850
rect 118130 82798 118132 82850
rect 118076 82404 118132 82798
rect 118076 82338 118132 82348
rect 117964 79940 118020 79950
rect 117964 79826 118020 79884
rect 117964 79774 117966 79826
rect 118018 79774 118020 79826
rect 117964 79762 118020 79774
rect 117964 78596 118020 78606
rect 117964 78258 118020 78540
rect 117964 78206 117966 78258
rect 118018 78206 118020 78258
rect 117964 78194 118020 78206
rect 118076 78594 118132 78606
rect 118076 78542 118078 78594
rect 118130 78542 118132 78594
rect 118076 78148 118132 78542
rect 118076 78082 118132 78092
rect 118076 70756 118132 70766
rect 118076 70662 118132 70700
rect 117068 57922 117124 57932
rect 117180 57932 117572 57988
rect 117628 67172 117796 67228
rect 117628 64932 117684 67172
rect 117964 67058 118020 67070
rect 117964 67006 117966 67058
rect 118018 67006 118020 67058
rect 117964 66948 118020 67006
rect 117964 66882 118020 66892
rect 117740 66276 117796 66286
rect 117740 65492 117796 66220
rect 117852 66164 117908 66174
rect 117852 66070 117908 66108
rect 117852 65492 117908 65502
rect 117740 65490 117908 65492
rect 117740 65438 117854 65490
rect 117906 65438 117908 65490
rect 117740 65436 117908 65438
rect 117852 65426 117908 65436
rect 117068 57764 117124 57774
rect 117180 57764 117236 57932
rect 117068 57762 117236 57764
rect 117068 57710 117070 57762
rect 117122 57710 117236 57762
rect 117068 57708 117236 57710
rect 117068 57698 117124 57708
rect 117292 57650 117348 57662
rect 117292 57598 117294 57650
rect 117346 57598 117348 57650
rect 116508 57540 116564 57550
rect 117292 57540 117348 57598
rect 116508 57538 117348 57540
rect 116508 57486 116510 57538
rect 116562 57486 117348 57538
rect 116508 57484 117348 57486
rect 115836 55972 115892 55982
rect 115836 55878 115892 55916
rect 116508 55468 116564 57484
rect 117628 55468 117684 64876
rect 118076 56644 118132 56654
rect 118076 56550 118132 56588
rect 115836 55410 115892 55422
rect 115836 55358 115838 55410
rect 115890 55358 115892 55410
rect 115836 54628 115892 55358
rect 115836 54562 115892 54572
rect 116060 55412 116564 55468
rect 117292 55412 117684 55468
rect 115500 50706 115556 50718
rect 115500 50654 115502 50706
rect 115554 50654 115556 50706
rect 115500 49924 115556 50654
rect 115500 49858 115556 49868
rect 115500 49138 115556 49150
rect 115500 49086 115502 49138
rect 115554 49086 115556 49138
rect 115500 48580 115556 49086
rect 115500 48514 115556 48524
rect 115500 48130 115556 48142
rect 115500 48078 115502 48130
rect 115554 48078 115556 48130
rect 115500 47908 115556 48078
rect 115500 47842 115556 47852
rect 115164 44884 115220 44894
rect 114940 43428 114996 43438
rect 114940 43334 114996 43372
rect 114380 41972 114436 41982
rect 114380 41878 114436 41916
rect 114940 41972 114996 41982
rect 114940 41878 114996 41916
rect 115164 40290 115220 44828
rect 115388 44548 115444 45276
rect 115500 46002 115556 46014
rect 115500 45950 115502 46002
rect 115554 45950 115556 46002
rect 115500 45220 115556 45950
rect 115500 45154 115556 45164
rect 115388 44482 115444 44492
rect 115836 41860 115892 41870
rect 115836 41766 115892 41804
rect 115500 41298 115556 41310
rect 115500 41246 115502 41298
rect 115554 41246 115556 41298
rect 115164 40238 115166 40290
rect 115218 40238 115220 40290
rect 115164 40226 115220 40238
rect 115276 41188 115332 41198
rect 114828 37828 114884 37838
rect 114828 36594 114884 37772
rect 114828 36542 114830 36594
rect 114882 36542 114884 36594
rect 114828 36530 114884 36542
rect 114492 35700 114548 35710
rect 114492 35606 114548 35644
rect 114940 35700 114996 35710
rect 114940 35606 114996 35644
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 112588 32340 112644 33516
rect 112588 32274 112644 32284
rect 112812 35252 112868 35262
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 110012 21522 110068 21532
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 112364 17668 112420 17678
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 111996 14074 112260 14084
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 112364 6130 112420 17612
rect 112364 6078 112366 6130
rect 112418 6078 112420 6130
rect 112364 5908 112420 6078
rect 112364 5842 112420 5852
rect 112812 5234 112868 35196
rect 115164 34130 115220 34142
rect 115164 34078 115166 34130
rect 115218 34078 115220 34130
rect 114604 34020 114660 34030
rect 114604 33926 114660 33964
rect 115164 34020 115220 34078
rect 115164 33954 115220 33964
rect 114940 32676 114996 32686
rect 114940 32582 114996 32620
rect 115276 31948 115332 41132
rect 115500 40516 115556 41246
rect 115500 40450 115556 40460
rect 116060 40180 116116 55412
rect 116284 53058 116340 53070
rect 116284 53006 116286 53058
rect 116338 53006 116340 53058
rect 116284 52612 116340 53006
rect 116284 52546 116340 52556
rect 116844 52834 116900 52846
rect 116844 52782 116846 52834
rect 116898 52782 116900 52834
rect 116844 52612 116900 52782
rect 116844 52546 116900 52556
rect 116172 50596 116228 50606
rect 116172 50594 117124 50596
rect 116172 50542 116174 50594
rect 116226 50542 117124 50594
rect 116172 50540 117124 50542
rect 116172 50530 116228 50540
rect 117068 50482 117124 50540
rect 117068 50430 117070 50482
rect 117122 50430 117124 50482
rect 117068 50418 117124 50430
rect 117292 50594 117348 55412
rect 117292 50542 117294 50594
rect 117346 50542 117348 50594
rect 116844 50036 116900 50046
rect 117292 50036 117348 50542
rect 116844 50034 117348 50036
rect 116844 49982 116846 50034
rect 116898 49982 117348 50034
rect 116844 49980 117348 49982
rect 116844 49970 116900 49980
rect 116172 49028 116228 49038
rect 116172 49026 117124 49028
rect 116172 48974 116174 49026
rect 116226 48974 117124 49026
rect 116172 48972 117124 48974
rect 116172 48962 116228 48972
rect 116956 48804 117012 48814
rect 116956 48710 117012 48748
rect 117068 48466 117124 48972
rect 117068 48414 117070 48466
rect 117122 48414 117124 48466
rect 117068 48402 117124 48414
rect 117292 48804 117348 48814
rect 116172 48244 116228 48254
rect 116172 48242 117124 48244
rect 116172 48190 116174 48242
rect 116226 48190 117124 48242
rect 116172 48188 117124 48190
rect 116172 48178 116228 48188
rect 117068 47346 117124 48188
rect 117068 47294 117070 47346
rect 117122 47294 117124 47346
rect 117068 47282 117124 47294
rect 117292 48242 117348 48748
rect 117292 48190 117294 48242
rect 117346 48190 117348 48242
rect 117292 47458 117348 48190
rect 117292 47406 117294 47458
rect 117346 47406 117348 47458
rect 116284 47234 116340 47246
rect 116284 47182 116286 47234
rect 116338 47182 116340 47234
rect 116284 47124 116340 47182
rect 117292 47124 117348 47406
rect 116284 47068 117348 47124
rect 116172 45892 116228 45902
rect 116172 45890 117124 45892
rect 116172 45838 116174 45890
rect 116226 45838 117124 45890
rect 116172 45836 117124 45838
rect 116172 45826 116228 45836
rect 116508 45332 116564 45342
rect 116508 45238 116564 45276
rect 117068 45330 117124 45836
rect 117068 45278 117070 45330
rect 117122 45278 117124 45330
rect 117068 45266 117124 45278
rect 116284 43650 116340 43662
rect 116284 43598 116286 43650
rect 116338 43598 116340 43650
rect 116284 43204 116340 43598
rect 116284 43138 116340 43148
rect 116844 43426 116900 43438
rect 116844 43374 116846 43426
rect 116898 43374 116900 43426
rect 116844 43204 116900 43374
rect 116844 43138 116900 43148
rect 116172 41188 116228 41198
rect 116172 41186 117124 41188
rect 116172 41134 116174 41186
rect 116226 41134 117124 41186
rect 116172 41132 117124 41134
rect 116172 41122 116228 41132
rect 116956 40962 117012 40974
rect 116956 40910 116958 40962
rect 117010 40910 117012 40962
rect 116060 40114 116116 40124
rect 116284 40514 116340 40526
rect 116284 40462 116286 40514
rect 116338 40462 116340 40514
rect 116284 39732 116340 40462
rect 116956 40404 117012 40910
rect 117068 40626 117124 41132
rect 117068 40574 117070 40626
rect 117122 40574 117124 40626
rect 117068 40562 117124 40574
rect 117292 40404 117348 47068
rect 118076 46786 118132 46798
rect 118076 46734 118078 46786
rect 118130 46734 118132 46786
rect 118076 46564 118132 46734
rect 118076 46498 118132 46508
rect 117404 45332 117460 45342
rect 117404 45218 117460 45276
rect 117404 45166 117406 45218
rect 117458 45166 117460 45218
rect 117404 45154 117460 45166
rect 118188 43764 118244 116508
rect 118300 115220 118356 119200
rect 118300 115154 118356 115164
rect 118188 43698 118244 43708
rect 116956 40402 117348 40404
rect 116956 40350 117294 40402
rect 117346 40350 117348 40402
rect 116956 40348 117348 40350
rect 116284 39666 116340 39676
rect 117068 39732 117124 39742
rect 117068 39638 117124 39676
rect 115612 39284 115668 39294
rect 115500 33684 115556 33694
rect 115500 33458 115556 33628
rect 115500 33406 115502 33458
rect 115554 33406 115556 33458
rect 115500 33394 115556 33406
rect 115388 32450 115444 32462
rect 115388 32398 115390 32450
rect 115442 32398 115444 32450
rect 115388 32340 115444 32398
rect 115388 32274 115444 32284
rect 115164 31892 115332 31948
rect 114380 30212 114436 30222
rect 114380 30118 114436 30156
rect 114940 30210 114996 30222
rect 114940 30158 114942 30210
rect 114994 30158 114996 30210
rect 114940 29988 114996 30158
rect 114940 29922 114996 29932
rect 114380 26292 114436 26302
rect 114380 26198 114436 26236
rect 114940 26292 114996 26302
rect 114940 26198 114996 26236
rect 114716 24500 114772 24510
rect 114492 15428 114548 15438
rect 114492 15334 114548 15372
rect 114492 14532 114548 14542
rect 114492 14438 114548 14476
rect 114492 8260 114548 8270
rect 114492 8166 114548 8204
rect 113148 5908 113204 5918
rect 113148 5814 113204 5852
rect 113820 5796 113876 5806
rect 112812 5182 112814 5234
rect 112866 5182 112868 5234
rect 112812 5170 112868 5182
rect 113708 5794 113876 5796
rect 113708 5742 113822 5794
rect 113874 5742 113876 5794
rect 113708 5740 113876 5742
rect 111356 5012 111412 5022
rect 111356 4918 111412 4956
rect 111916 5012 111972 5022
rect 111916 4918 111972 4956
rect 112252 4900 112308 4938
rect 112252 4834 112308 4844
rect 113148 4900 113204 4910
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 111996 4666 112260 4676
rect 112364 4340 112420 4350
rect 112364 4246 112420 4284
rect 113148 4338 113204 4844
rect 113148 4286 113150 4338
rect 113202 4286 113204 4338
rect 113148 4274 113204 4286
rect 111692 4228 111748 4238
rect 111692 4134 111748 4172
rect 108332 3602 108388 3612
rect 111580 3668 111636 3678
rect 111580 3574 111636 3612
rect 103852 3502 103854 3554
rect 103906 3502 103908 3554
rect 103852 3490 103908 3502
rect 112364 3556 112420 3566
rect 110908 3444 110964 3454
rect 105532 3330 105588 3342
rect 109116 3332 109172 3342
rect 109788 3332 109844 3342
rect 105532 3278 105534 3330
rect 105586 3278 105588 3330
rect 104300 1762 104356 1774
rect 104300 1710 104302 1762
rect 104354 1710 104356 1762
rect 104300 800 104356 1710
rect 105532 1762 105588 3278
rect 105532 1710 105534 1762
rect 105586 1710 105588 1762
rect 105532 1698 105588 1710
rect 109004 3330 109172 3332
rect 109004 3278 109118 3330
rect 109170 3278 109172 3330
rect 109004 3276 109172 3278
rect 109004 800 109060 3276
rect 109116 3266 109172 3276
rect 109676 3330 109844 3332
rect 109676 3278 109790 3330
rect 109842 3278 109844 3330
rect 109676 3276 109844 3278
rect 109676 800 109732 3276
rect 109788 3266 109844 3276
rect 110908 800 110964 3388
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 112364 800 112420 3500
rect 112588 3444 112644 3454
rect 112588 3350 112644 3388
rect 113708 800 113764 5740
rect 113820 5730 113876 5740
rect 114716 5236 114772 24444
rect 115164 21028 115220 31892
rect 115500 30882 115556 30894
rect 115500 30830 115502 30882
rect 115554 30830 115556 30882
rect 115500 30436 115556 30830
rect 115500 30370 115556 30380
rect 115500 30212 115556 30222
rect 115612 30212 115668 39228
rect 117292 39284 117348 40348
rect 117292 39218 117348 39228
rect 118076 38946 118132 38958
rect 118076 38894 118078 38946
rect 118130 38894 118132 38946
rect 118076 38724 118132 38894
rect 118076 38658 118132 38668
rect 116172 36372 116228 36382
rect 116172 36278 116228 36316
rect 117068 36372 117124 36382
rect 117068 36258 117124 36316
rect 117068 36206 117070 36258
rect 117122 36206 117124 36258
rect 117068 35812 117124 36206
rect 117068 35746 117124 35756
rect 115836 35586 115892 35598
rect 115836 35534 115838 35586
rect 115890 35534 115892 35586
rect 115836 35140 115892 35534
rect 115836 35074 115892 35084
rect 116172 34914 116228 34926
rect 116172 34862 116174 34914
rect 116226 34862 116228 34914
rect 115948 34690 116004 34702
rect 115948 34638 115950 34690
rect 116002 34638 116004 34690
rect 115948 34242 116004 34638
rect 115948 34190 115950 34242
rect 116002 34190 116004 34242
rect 115948 34178 116004 34190
rect 116060 34020 116116 34030
rect 116060 33346 116116 33964
rect 116060 33294 116062 33346
rect 116114 33294 116116 33346
rect 116060 33282 116116 33294
rect 116060 32788 116116 32798
rect 116172 32788 116228 34862
rect 116060 32786 116228 32788
rect 116060 32734 116062 32786
rect 116114 32734 116228 32786
rect 116060 32732 116228 32734
rect 117180 34020 117236 34030
rect 116060 32722 116116 32732
rect 116620 32676 116676 32686
rect 116620 32582 116676 32620
rect 117180 32674 117236 33964
rect 118076 34020 118132 34030
rect 118076 33926 118132 33964
rect 117180 32622 117182 32674
rect 117234 32622 117236 32674
rect 117180 32610 117236 32622
rect 116396 32340 116452 32350
rect 116172 30994 116228 31006
rect 116172 30942 116174 30994
rect 116226 30942 116228 30994
rect 116172 30434 116228 30942
rect 116172 30382 116174 30434
rect 116226 30382 116228 30434
rect 116172 30370 116228 30382
rect 115556 30156 115668 30212
rect 115500 30080 115556 30156
rect 116284 29988 116340 29998
rect 116284 29894 116340 29932
rect 115500 27186 115556 27198
rect 115500 27134 115502 27186
rect 115554 27134 115556 27186
rect 115500 27076 115556 27134
rect 115500 27010 115556 27020
rect 116172 27074 116228 27086
rect 116172 27022 116174 27074
rect 116226 27022 116228 27074
rect 116172 26964 116228 27022
rect 116172 26898 116228 26908
rect 115836 26178 115892 26190
rect 115836 26126 115838 26178
rect 115890 26126 115892 26178
rect 115836 25732 115892 26126
rect 116396 26068 116452 32284
rect 116508 30436 116564 30446
rect 116508 30434 117124 30436
rect 116508 30382 116510 30434
rect 116562 30382 117124 30434
rect 116508 30380 117124 30382
rect 116508 30370 116564 30380
rect 117068 30098 117124 30380
rect 117068 30046 117070 30098
rect 117122 30046 117124 30098
rect 117068 30034 117124 30046
rect 117404 30098 117460 30110
rect 117404 30046 117406 30098
rect 117458 30046 117460 30098
rect 117404 29988 117460 30046
rect 117068 26964 117124 26974
rect 117068 26870 117124 26908
rect 117404 26962 117460 29932
rect 117404 26910 117406 26962
rect 117458 26910 117460 26962
rect 116732 26516 116788 26526
rect 117404 26516 117460 26910
rect 116732 26514 117460 26516
rect 116732 26462 116734 26514
rect 116786 26462 117460 26514
rect 116732 26460 117460 26462
rect 116732 26450 116788 26460
rect 116396 26012 116676 26068
rect 115836 25666 115892 25676
rect 116620 23492 116676 26012
rect 116620 23436 117348 23492
rect 116620 23378 116676 23436
rect 116620 23326 116622 23378
rect 116674 23326 116676 23378
rect 116620 23314 116676 23326
rect 117068 23266 117124 23278
rect 117068 23214 117070 23266
rect 117122 23214 117124 23266
rect 115500 22482 115556 22494
rect 115500 22430 115502 22482
rect 115554 22430 115556 22482
rect 115500 22372 115556 22430
rect 115500 22306 115556 22316
rect 116172 22372 116228 22382
rect 117068 22372 117124 23214
rect 117292 23154 117348 23436
rect 117292 23102 117294 23154
rect 117346 23102 117348 23154
rect 117292 23090 117348 23102
rect 116172 22370 117124 22372
rect 116172 22318 116174 22370
rect 116226 22318 117124 22370
rect 116172 22316 117124 22318
rect 116172 22306 116228 22316
rect 115164 20962 115220 20972
rect 115500 19346 115556 19358
rect 115500 19294 115502 19346
rect 115554 19294 115556 19346
rect 115500 19012 115556 19294
rect 116172 19236 116228 19246
rect 117404 19236 117460 26460
rect 116172 19234 117124 19236
rect 116172 19182 116174 19234
rect 116226 19182 117124 19234
rect 116172 19180 117124 19182
rect 116172 19170 116228 19180
rect 117068 19122 117124 19180
rect 117068 19070 117070 19122
rect 117122 19070 117124 19122
rect 117068 19058 117124 19070
rect 117180 19234 117460 19236
rect 117180 19182 117406 19234
rect 117458 19182 117460 19234
rect 117180 19180 117460 19182
rect 115500 18946 115556 18956
rect 117180 18788 117236 19180
rect 117404 19170 117460 19180
rect 116732 18732 117236 18788
rect 116732 18674 116788 18732
rect 116732 18622 116734 18674
rect 116786 18622 116788 18674
rect 116732 18610 116788 18622
rect 114940 15428 114996 15438
rect 114940 15314 114996 15372
rect 114940 15262 114942 15314
rect 114994 15262 114996 15314
rect 114940 15250 114996 15262
rect 115836 15202 115892 15214
rect 115836 15150 115838 15202
rect 115890 15150 115892 15202
rect 115836 14980 115892 15150
rect 115836 14914 115892 14924
rect 115836 14642 115892 14654
rect 115836 14590 115838 14642
rect 115890 14590 115892 14642
rect 114940 14532 114996 14542
rect 114940 14438 114996 14476
rect 115836 14308 115892 14590
rect 115836 14242 115892 14252
rect 116284 12290 116340 12302
rect 116284 12238 116286 12290
rect 116338 12238 116340 12290
rect 114940 12068 114996 12078
rect 114940 11974 114996 12012
rect 116284 11844 116340 12238
rect 116284 11778 116340 11788
rect 116844 12066 116900 12078
rect 116844 12014 116846 12066
rect 116898 12014 116900 12066
rect 116844 11844 116900 12014
rect 116844 11778 116900 11788
rect 115500 9938 115556 9950
rect 115500 9886 115502 9938
rect 115554 9886 115556 9938
rect 115500 9604 115556 9886
rect 116172 9828 116228 9838
rect 117180 9828 117236 18732
rect 118076 16996 118132 17006
rect 118076 16902 118132 16940
rect 117292 9828 117348 9838
rect 116172 9826 117124 9828
rect 116172 9774 116174 9826
rect 116226 9774 117124 9826
rect 116172 9772 117124 9774
rect 116172 9762 116228 9772
rect 117068 9714 117124 9772
rect 117068 9662 117070 9714
rect 117122 9662 117124 9714
rect 117068 9650 117124 9662
rect 117180 9826 117348 9828
rect 117180 9774 117294 9826
rect 117346 9774 117348 9826
rect 117180 9772 117348 9774
rect 115500 9538 115556 9548
rect 117180 9492 117236 9772
rect 116732 9436 117236 9492
rect 116732 9266 116788 9436
rect 116732 9214 116734 9266
rect 116786 9214 116788 9266
rect 116732 9202 116788 9214
rect 117292 8428 117348 9772
rect 115836 8370 115892 8382
rect 117292 8372 117460 8428
rect 115836 8318 115838 8370
rect 115890 8318 115892 8370
rect 114940 8260 114996 8270
rect 114940 8166 114996 8204
rect 115836 8260 115892 8318
rect 115836 8194 115892 8204
rect 116620 7532 117124 7588
rect 116172 7476 116228 7486
rect 116620 7476 116676 7532
rect 116172 7474 116676 7476
rect 116172 7422 116174 7474
rect 116226 7422 116676 7474
rect 116172 7420 116676 7422
rect 116172 7410 116228 7420
rect 115500 7362 115556 7374
rect 115500 7310 115502 7362
rect 115554 7310 115556 7362
rect 115500 6916 115556 7310
rect 115500 6850 115556 6860
rect 116732 7362 116788 7374
rect 116732 7310 116734 7362
rect 116786 7310 116788 7362
rect 114828 6804 114884 6814
rect 114828 6710 114884 6748
rect 116172 6578 116228 6590
rect 116172 6526 116174 6578
rect 116226 6526 116228 6578
rect 116172 6244 116228 6526
rect 116172 6178 116228 6188
rect 116732 6244 116788 7310
rect 117068 6578 117124 7532
rect 117068 6526 117070 6578
rect 117122 6526 117124 6578
rect 117068 6514 117124 6526
rect 117404 6578 117460 8372
rect 117404 6526 117406 6578
rect 117458 6526 117460 6578
rect 116732 6178 116788 6188
rect 114940 6020 114996 6030
rect 114940 5794 114996 5964
rect 116284 6018 116340 6030
rect 116284 5966 116286 6018
rect 116338 5966 116340 6018
rect 114940 5742 114942 5794
rect 114994 5742 114996 5794
rect 114940 5730 114996 5742
rect 115500 5796 115556 5806
rect 114828 5236 114884 5246
rect 114716 5234 114884 5236
rect 114716 5182 114830 5234
rect 114882 5182 114884 5234
rect 114716 5180 114884 5182
rect 114828 5170 114884 5180
rect 114156 5012 114212 5022
rect 114156 5010 114548 5012
rect 114156 4958 114158 5010
rect 114210 4958 114548 5010
rect 114156 4956 114548 4958
rect 114156 4946 114212 4956
rect 113820 4226 113876 4238
rect 113820 4174 113822 4226
rect 113874 4174 113876 4226
rect 113820 3556 113876 4174
rect 113820 3490 113876 3500
rect 114156 3444 114212 3454
rect 114268 3444 114324 3454
rect 114156 3442 114268 3444
rect 114156 3390 114158 3442
rect 114210 3390 114268 3442
rect 114156 3388 114268 3390
rect 114156 3378 114212 3388
rect 114268 800 114324 3388
rect 114492 3442 114548 4956
rect 114940 4452 114996 4462
rect 114940 4226 114996 4396
rect 114940 4174 114942 4226
rect 114994 4174 114996 4226
rect 114940 4162 114996 4174
rect 115500 3666 115556 5740
rect 116172 5010 116228 5022
rect 116172 4958 116174 5010
rect 116226 4958 116228 5010
rect 116172 4900 116228 4958
rect 116284 5012 116340 5966
rect 116284 4946 116340 4956
rect 116844 5794 116900 5806
rect 116844 5742 116846 5794
rect 116898 5742 116900 5794
rect 116172 4834 116228 4844
rect 116844 4788 116900 5742
rect 117292 5794 117348 5806
rect 117292 5742 117294 5794
rect 117346 5742 117348 5794
rect 117292 5012 117348 5742
rect 117068 4900 117124 4910
rect 117068 4806 117124 4844
rect 116844 4722 116900 4732
rect 117292 4564 117348 4956
rect 117292 4498 117348 4508
rect 117404 4788 117460 6526
rect 116284 4452 116340 4462
rect 116284 4358 116340 4396
rect 117068 4450 117124 4462
rect 117068 4398 117070 4450
rect 117122 4398 117124 4450
rect 117068 4340 117124 4398
rect 117068 4274 117124 4284
rect 117404 4450 117460 4732
rect 118860 4564 118916 4574
rect 117404 4398 117406 4450
rect 117458 4398 117460 4450
rect 115500 3614 115502 3666
rect 115554 3614 115556 3666
rect 115500 3602 115556 3614
rect 117404 3666 117460 4398
rect 117852 4452 117908 4462
rect 117404 3614 117406 3666
rect 117458 3614 117460 3666
rect 117404 3602 117460 3614
rect 117628 4228 117684 4238
rect 114492 3390 114494 3442
rect 114546 3390 114548 3442
rect 114492 1540 114548 3390
rect 116508 3444 116564 3454
rect 116508 3350 116564 3388
rect 114492 1474 114548 1484
rect 117628 800 117684 4172
rect 117852 4226 117908 4396
rect 117852 4174 117854 4226
rect 117906 4174 117908 4226
rect 117852 3556 117908 4174
rect 117852 3490 117908 3500
rect 118076 3330 118132 3342
rect 118076 3278 118078 3330
rect 118130 3278 118132 3330
rect 118076 2212 118132 3278
rect 118076 2146 118132 2156
rect 118860 800 118916 4508
rect 100744 200 100968 728
rect 101416 200 101640 728
rect 101724 700 102452 756
rect 102760 728 103012 800
rect 104104 728 104356 800
rect 102760 200 102984 728
rect 104104 200 104328 728
rect 105448 200 105672 800
rect 106120 200 106344 800
rect 107464 200 107688 800
rect 108808 728 109060 800
rect 109480 728 109732 800
rect 108808 200 109032 728
rect 109480 200 109704 728
rect 110824 200 111048 800
rect 112168 728 112420 800
rect 113512 728 113764 800
rect 112168 200 112392 728
rect 113512 200 113736 728
rect 114184 200 114408 800
rect 115528 200 115752 800
rect 116872 200 117096 800
rect 117544 200 117768 800
rect 118860 728 119112 800
rect 118888 200 119112 728
<< via2 >>
rect 140 117852 196 117908
rect 2044 118860 2100 118916
rect 1820 117852 1876 117908
rect 1932 115948 1988 116004
rect 3388 116620 3444 116676
rect 3052 116172 3108 116228
rect 4476 116842 4532 116844
rect 4476 116790 4478 116842
rect 4478 116790 4530 116842
rect 4530 116790 4532 116842
rect 4476 116788 4532 116790
rect 4580 116842 4636 116844
rect 4580 116790 4582 116842
rect 4582 116790 4634 116842
rect 4634 116790 4636 116842
rect 4580 116788 4636 116790
rect 4684 116842 4740 116844
rect 4684 116790 4686 116842
rect 4686 116790 4738 116842
rect 4738 116790 4740 116842
rect 4684 116788 4740 116790
rect 3836 116226 3892 116228
rect 3836 116174 3838 116226
rect 3838 116174 3890 116226
rect 3890 116174 3892 116226
rect 3836 116172 3892 116174
rect 5740 115890 5796 115892
rect 5740 115838 5742 115890
rect 5742 115838 5794 115890
rect 5794 115838 5796 115890
rect 5740 115836 5796 115838
rect 4732 115724 4788 115780
rect 3164 114940 3220 114996
rect 3052 114882 3108 114884
rect 3052 114830 3054 114882
rect 3054 114830 3106 114882
rect 3106 114830 3108 114882
rect 3052 114828 3108 114830
rect 2380 114604 2436 114660
rect 1820 113484 1876 113540
rect 1932 112418 1988 112420
rect 1932 112366 1934 112418
rect 1934 112366 1986 112418
rect 1986 112366 1988 112418
rect 1932 112364 1988 112366
rect 1708 111074 1764 111076
rect 1708 111022 1710 111074
rect 1710 111022 1762 111074
rect 1762 111022 1764 111074
rect 1708 111020 1764 111022
rect 1820 109676 1876 109732
rect 1820 107660 1876 107716
rect 1932 104300 1988 104356
rect 1932 103010 1988 103012
rect 1932 102958 1934 103010
rect 1934 102958 1986 103010
rect 1986 102958 1988 103010
rect 1932 102956 1988 102958
rect 3612 114940 3668 114996
rect 3836 114940 3892 114996
rect 3724 114828 3780 114884
rect 5292 115554 5348 115556
rect 5292 115502 5294 115554
rect 5294 115502 5346 115554
rect 5346 115502 5348 115554
rect 5292 115500 5348 115502
rect 4476 115274 4532 115276
rect 4476 115222 4478 115274
rect 4478 115222 4530 115274
rect 4530 115222 4532 115274
rect 4476 115220 4532 115222
rect 4580 115274 4636 115276
rect 4580 115222 4582 115274
rect 4582 115222 4634 115274
rect 4634 115222 4636 115274
rect 4580 115220 4636 115222
rect 4684 115274 4740 115276
rect 4684 115222 4686 115274
rect 4686 115222 4738 115274
rect 4738 115222 4740 115274
rect 4684 115220 4740 115222
rect 4396 114994 4452 114996
rect 4396 114942 4398 114994
rect 4398 114942 4450 114994
rect 4450 114942 4452 114994
rect 4396 114940 4452 114942
rect 5292 114940 5348 114996
rect 3724 113932 3780 113988
rect 3388 113820 3444 113876
rect 4476 113706 4532 113708
rect 4476 113654 4478 113706
rect 4478 113654 4530 113706
rect 4530 113654 4532 113706
rect 4476 113652 4532 113654
rect 4580 113706 4636 113708
rect 4580 113654 4582 113706
rect 4582 113654 4634 113706
rect 4634 113654 4636 113706
rect 4580 113652 4636 113654
rect 4684 113706 4740 113708
rect 4684 113654 4686 113706
rect 4686 113654 4738 113706
rect 4738 113654 4740 113706
rect 4684 113652 4740 113654
rect 2380 101666 2436 101668
rect 2380 101614 2382 101666
rect 2382 101614 2434 101666
rect 2434 101614 2436 101666
rect 2380 101612 2436 101614
rect 1820 100940 1876 100996
rect 1820 99372 1876 99428
rect 2604 99202 2660 99204
rect 2604 99150 2606 99202
rect 2606 99150 2658 99202
rect 2658 99150 2660 99202
rect 2604 99148 2660 99150
rect 1932 98306 1988 98308
rect 1932 98254 1934 98306
rect 1934 98254 1986 98306
rect 1986 98254 1988 98306
rect 1932 98252 1988 98254
rect 1708 96962 1764 96964
rect 1708 96910 1710 96962
rect 1710 96910 1762 96962
rect 1762 96910 1764 96962
rect 1708 96908 1764 96910
rect 1932 94892 1988 94948
rect 4476 112138 4532 112140
rect 4476 112086 4478 112138
rect 4478 112086 4530 112138
rect 4530 112086 4532 112138
rect 4476 112084 4532 112086
rect 4580 112138 4636 112140
rect 4580 112086 4582 112138
rect 4582 112086 4634 112138
rect 4634 112086 4636 112138
rect 4580 112084 4636 112086
rect 4684 112138 4740 112140
rect 4684 112086 4686 112138
rect 4686 112086 4738 112138
rect 4738 112086 4740 112138
rect 4684 112084 4740 112086
rect 3276 111858 3332 111860
rect 3276 111806 3278 111858
rect 3278 111806 3330 111858
rect 3330 111806 3332 111858
rect 3276 111804 3332 111806
rect 4476 110570 4532 110572
rect 4476 110518 4478 110570
rect 4478 110518 4530 110570
rect 4530 110518 4532 110570
rect 4476 110516 4532 110518
rect 4580 110570 4636 110572
rect 4580 110518 4582 110570
rect 4582 110518 4634 110570
rect 4634 110518 4636 110570
rect 4580 110516 4636 110518
rect 4684 110570 4740 110572
rect 4684 110518 4686 110570
rect 4686 110518 4738 110570
rect 4738 110518 4740 110570
rect 4684 110516 4740 110518
rect 4476 109002 4532 109004
rect 4476 108950 4478 109002
rect 4478 108950 4530 109002
rect 4530 108950 4532 109002
rect 4476 108948 4532 108950
rect 4580 109002 4636 109004
rect 4580 108950 4582 109002
rect 4582 108950 4634 109002
rect 4634 108950 4636 109002
rect 4580 108948 4636 108950
rect 4684 109002 4740 109004
rect 4684 108950 4686 109002
rect 4686 108950 4738 109002
rect 4738 108950 4740 109002
rect 4684 108948 4740 108950
rect 4476 107434 4532 107436
rect 4476 107382 4478 107434
rect 4478 107382 4530 107434
rect 4530 107382 4532 107434
rect 4476 107380 4532 107382
rect 4580 107434 4636 107436
rect 4580 107382 4582 107434
rect 4582 107382 4634 107434
rect 4634 107382 4636 107434
rect 4580 107380 4636 107382
rect 4684 107434 4740 107436
rect 4684 107382 4686 107434
rect 4686 107382 4738 107434
rect 4738 107382 4740 107434
rect 4684 107380 4740 107382
rect 4476 105866 4532 105868
rect 4476 105814 4478 105866
rect 4478 105814 4530 105866
rect 4530 105814 4532 105866
rect 4476 105812 4532 105814
rect 4580 105866 4636 105868
rect 4580 105814 4582 105866
rect 4582 105814 4634 105866
rect 4634 105814 4636 105866
rect 4580 105812 4636 105814
rect 4684 105866 4740 105868
rect 4684 105814 4686 105866
rect 4686 105814 4738 105866
rect 4738 105814 4740 105866
rect 4684 105812 4740 105814
rect 3052 104524 3108 104580
rect 3612 104578 3668 104580
rect 3612 104526 3614 104578
rect 3614 104526 3666 104578
rect 3666 104526 3668 104578
rect 3612 104524 3668 104526
rect 4476 104298 4532 104300
rect 4476 104246 4478 104298
rect 4478 104246 4530 104298
rect 4530 104246 4532 104298
rect 4476 104244 4532 104246
rect 4580 104298 4636 104300
rect 4580 104246 4582 104298
rect 4582 104246 4634 104298
rect 4634 104246 4636 104298
rect 4580 104244 4636 104246
rect 4684 104298 4740 104300
rect 4684 104246 4686 104298
rect 4686 104246 4738 104298
rect 4738 104246 4740 104298
rect 4684 104244 4740 104246
rect 3052 102956 3108 103012
rect 3612 103010 3668 103012
rect 3612 102958 3614 103010
rect 3614 102958 3666 103010
rect 3666 102958 3668 103010
rect 3612 102956 3668 102958
rect 4476 102730 4532 102732
rect 4476 102678 4478 102730
rect 4478 102678 4530 102730
rect 4530 102678 4532 102730
rect 4476 102676 4532 102678
rect 4580 102730 4636 102732
rect 4580 102678 4582 102730
rect 4582 102678 4634 102730
rect 4634 102678 4636 102730
rect 4580 102676 4636 102678
rect 4684 102730 4740 102732
rect 4684 102678 4686 102730
rect 4686 102678 4738 102730
rect 4738 102678 4740 102730
rect 4684 102676 4740 102678
rect 3164 102450 3220 102452
rect 3164 102398 3166 102450
rect 3166 102398 3218 102450
rect 3218 102398 3220 102450
rect 3164 102396 3220 102398
rect 4476 101162 4532 101164
rect 4476 101110 4478 101162
rect 4478 101110 4530 101162
rect 4530 101110 4532 101162
rect 4476 101108 4532 101110
rect 4580 101162 4636 101164
rect 4580 101110 4582 101162
rect 4582 101110 4634 101162
rect 4634 101110 4636 101162
rect 4580 101108 4636 101110
rect 4684 101162 4740 101164
rect 4684 101110 4686 101162
rect 4686 101110 4738 101162
rect 4738 101110 4740 101162
rect 4684 101108 4740 101110
rect 3276 99874 3332 99876
rect 3276 99822 3278 99874
rect 3278 99822 3330 99874
rect 3330 99822 3332 99874
rect 3276 99820 3332 99822
rect 4476 99594 4532 99596
rect 4476 99542 4478 99594
rect 4478 99542 4530 99594
rect 4530 99542 4532 99594
rect 4476 99540 4532 99542
rect 4580 99594 4636 99596
rect 4580 99542 4582 99594
rect 4582 99542 4634 99594
rect 4634 99542 4636 99594
rect 4580 99540 4636 99542
rect 4684 99594 4740 99596
rect 4684 99542 4686 99594
rect 4686 99542 4738 99594
rect 4738 99542 4740 99594
rect 4684 99540 4740 99542
rect 3164 99148 3220 99204
rect 4476 98026 4532 98028
rect 4476 97974 4478 98026
rect 4478 97974 4530 98026
rect 4530 97974 4532 98026
rect 4476 97972 4532 97974
rect 4580 98026 4636 98028
rect 4580 97974 4582 98026
rect 4582 97974 4634 98026
rect 4634 97974 4636 98026
rect 4580 97972 4636 97974
rect 4684 98026 4740 98028
rect 4684 97974 4686 98026
rect 4686 97974 4738 98026
rect 4738 97974 4740 98026
rect 4684 97972 4740 97974
rect 3276 97746 3332 97748
rect 3276 97694 3278 97746
rect 3278 97694 3330 97746
rect 3330 97694 3332 97746
rect 3276 97692 3332 97694
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 1932 93602 1988 93604
rect 1932 93550 1934 93602
rect 1934 93550 1986 93602
rect 1986 93550 1988 93602
rect 1932 93548 1988 93550
rect 1932 92818 1988 92820
rect 1932 92766 1934 92818
rect 1934 92766 1986 92818
rect 1986 92766 1988 92818
rect 1932 92764 1988 92766
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 3052 93548 3108 93604
rect 1932 90188 1988 90244
rect 1932 88898 1988 88900
rect 1932 88846 1934 88898
rect 1934 88846 1986 88898
rect 1986 88846 1988 88898
rect 1932 88844 1988 88846
rect 1932 88114 1988 88116
rect 1932 88062 1934 88114
rect 1934 88062 1986 88114
rect 1986 88062 1988 88114
rect 1932 88060 1988 88062
rect 1820 85484 1876 85540
rect 1820 84140 1876 84196
rect 1932 82124 1988 82180
rect 3052 89010 3108 89012
rect 3052 88958 3054 89010
rect 3054 88958 3106 89010
rect 3106 88958 3108 89010
rect 3052 88956 3108 88958
rect 1932 80108 1988 80164
rect 3612 93602 3668 93604
rect 3612 93550 3614 93602
rect 3614 93550 3666 93602
rect 3666 93550 3668 93602
rect 3612 93548 3668 93550
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 3276 93042 3332 93044
rect 3276 92990 3278 93042
rect 3278 92990 3330 93042
rect 3330 92990 3332 93042
rect 3276 92988 3332 92990
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 5068 89628 5124 89684
rect 3500 89010 3556 89012
rect 3500 88958 3502 89010
rect 3502 88958 3554 89010
rect 3554 88958 3556 89010
rect 3500 88956 3556 88958
rect 5068 88956 5124 89012
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 3276 88338 3332 88340
rect 3276 88286 3278 88338
rect 3278 88286 3330 88338
rect 3330 88286 3332 88338
rect 3276 88284 3332 88286
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 1932 78706 1988 78708
rect 1932 78654 1934 78706
rect 1934 78654 1986 78706
rect 1986 78654 1988 78706
rect 1932 78652 1988 78654
rect 1932 76076 1988 76132
rect 1932 75404 1988 75460
rect 2828 75010 2884 75012
rect 2828 74958 2830 75010
rect 2830 74958 2882 75010
rect 2882 74958 2884 75010
rect 2828 74956 2884 74958
rect 1820 71148 1876 71204
rect 2828 70364 2884 70420
rect 1932 69298 1988 69300
rect 1932 69246 1934 69298
rect 1934 69246 1986 69298
rect 1986 69246 1988 69298
rect 1932 69244 1988 69246
rect 1932 68012 1988 68068
rect 3052 78540 3108 78596
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 3500 78594 3556 78596
rect 3500 78542 3502 78594
rect 3502 78542 3554 78594
rect 3554 78542 3556 78594
rect 3500 78540 3556 78542
rect 5852 78540 5908 78596
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 4396 76242 4452 76244
rect 4396 76190 4398 76242
rect 4398 76190 4450 76242
rect 4450 76190 4452 76242
rect 4396 76188 4452 76190
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 3276 75122 3332 75124
rect 3276 75070 3278 75122
rect 3278 75070 3330 75122
rect 3330 75070 3332 75122
rect 3276 75068 3332 75070
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 3388 70924 3444 70980
rect 3388 70418 3444 70420
rect 3388 70366 3390 70418
rect 3390 70366 3442 70418
rect 3442 70366 3444 70418
rect 3388 70364 3444 70366
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 3052 68348 3108 68404
rect 3612 68348 3668 68404
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 1820 65772 1876 65828
rect 1932 63308 1988 63364
rect 1820 62578 1876 62580
rect 1820 62526 1822 62578
rect 1822 62526 1874 62578
rect 1874 62526 1876 62578
rect 1820 62524 1876 62526
rect 3052 61628 3108 61684
rect 1932 61292 1988 61348
rect 1932 59890 1988 59892
rect 1932 59838 1934 59890
rect 1934 59838 1986 59890
rect 1986 59838 1988 59890
rect 1932 59836 1988 59838
rect 1820 58546 1876 58548
rect 1820 58494 1822 58546
rect 1822 58494 1874 58546
rect 1874 58494 1876 58546
rect 1820 58492 1876 58494
rect 1932 56588 1988 56644
rect 3052 56588 3108 56644
rect 1820 54572 1876 54628
rect 1820 51660 1876 51716
rect 1820 48524 1876 48580
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 3276 66386 3332 66388
rect 3276 66334 3278 66386
rect 3278 66334 3330 66386
rect 3330 66334 3332 66386
rect 3276 66332 3332 66334
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 3388 64092 3444 64148
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 9772 115554 9828 115556
rect 9772 115502 9774 115554
rect 9774 115502 9826 115554
rect 9826 115502 9828 115554
rect 9772 115500 9828 115502
rect 10332 115500 10388 115556
rect 11340 115500 11396 115556
rect 11788 116562 11844 116564
rect 11788 116510 11790 116562
rect 11790 116510 11842 116562
rect 11842 116510 11844 116562
rect 11788 116508 11844 116510
rect 15708 116396 15764 116452
rect 12348 115612 12404 115668
rect 11900 114604 11956 114660
rect 7532 69692 7588 69748
rect 9212 113932 9268 113988
rect 3388 60172 3444 60228
rect 3276 59106 3332 59108
rect 3276 59054 3278 59106
rect 3278 59054 3330 59106
rect 3330 59054 3332 59106
rect 3276 59052 3332 59054
rect 5852 63196 5908 63252
rect 6748 68460 6804 68516
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 3612 61682 3668 61684
rect 3612 61630 3614 61682
rect 3614 61630 3666 61682
rect 3666 61630 3668 61682
rect 3612 61628 3668 61630
rect 6748 61628 6804 61684
rect 5852 60844 5908 60900
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 5852 60172 5908 60228
rect 5852 59388 5908 59444
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 3500 58156 3556 58212
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 3500 56642 3556 56644
rect 3500 56590 3502 56642
rect 3502 56590 3554 56642
rect 3554 56590 3556 56642
rect 3500 56588 3556 56590
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3388 51996 3444 52052
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 1932 46562 1988 46564
rect 1932 46510 1934 46562
rect 1934 46510 1986 46562
rect 1986 46510 1988 46562
rect 1932 46508 1988 46510
rect 3052 45612 3108 45668
rect 1932 45164 1988 45220
rect 1708 40514 1764 40516
rect 1708 40462 1710 40514
rect 1710 40462 1762 40514
rect 1762 40462 1764 40514
rect 1708 40460 1764 40462
rect 3052 39618 3108 39620
rect 3052 39566 3054 39618
rect 3054 39566 3106 39618
rect 3106 39566 3108 39618
rect 3052 39564 3108 39566
rect 1932 39116 1988 39172
rect 1932 37772 1988 37828
rect 3052 37772 3108 37828
rect 1932 37100 1988 37156
rect 2156 35810 2212 35812
rect 2156 35758 2158 35810
rect 2158 35758 2210 35810
rect 2210 35758 2212 35810
rect 2156 35756 2212 35758
rect 1932 34412 1988 34468
rect 3052 33964 3108 34020
rect 1932 33740 1988 33796
rect 1932 32172 1988 32228
rect 1820 29650 1876 29652
rect 1820 29598 1822 29650
rect 1822 29598 1874 29650
rect 1874 29598 1876 29650
rect 1820 29596 1876 29598
rect 1708 26402 1764 26404
rect 1708 26350 1710 26402
rect 1710 26350 1762 26402
rect 1762 26350 1764 26402
rect 1708 26348 1764 26350
rect 1932 25004 1988 25060
rect 3052 24556 3108 24612
rect 1932 24332 1988 24388
rect 1932 23042 1988 23044
rect 1932 22990 1934 23042
rect 1934 22990 1986 23042
rect 1986 22990 1988 23042
rect 1932 22988 1988 22990
rect 3052 22988 3108 23044
rect 1820 21420 1876 21476
rect 3052 21308 3108 21364
rect 1932 20972 1988 21028
rect 1820 18284 1876 18340
rect 1820 16940 1876 16996
rect 3052 16882 3108 16884
rect 3052 16830 3054 16882
rect 3054 16830 3106 16882
rect 3106 16830 3108 16882
rect 3052 16828 3108 16830
rect 1932 16268 1988 16324
rect 1932 11564 1988 11620
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3500 45666 3556 45668
rect 3500 45614 3502 45666
rect 3502 45614 3554 45666
rect 3554 45614 3556 45666
rect 3500 45612 3556 45614
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 3276 41298 3332 41300
rect 3276 41246 3278 41298
rect 3278 41246 3330 41298
rect 3330 41246 3332 41298
rect 3276 41244 3332 41246
rect 3612 41132 3668 41188
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3612 39564 3668 39620
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3388 37884 3444 37940
rect 3500 37826 3556 37828
rect 3500 37774 3502 37826
rect 3502 37774 3554 37826
rect 3554 37774 3556 37826
rect 3500 37772 3556 37774
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 3276 36594 3332 36596
rect 3276 36542 3278 36594
rect 3278 36542 3330 36594
rect 3330 36542 3332 36594
rect 3276 36540 3332 36542
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3388 35084 3444 35140
rect 3612 34018 3668 34020
rect 3612 33966 3614 34018
rect 3614 33966 3666 34018
rect 3666 33966 3668 34018
rect 3612 33964 3668 33966
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 3276 32450 3332 32452
rect 3276 32398 3278 32450
rect 3278 32398 3330 32450
rect 3330 32398 3332 32450
rect 3276 32396 3332 32398
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3388 30156 3444 30212
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3388 27244 3444 27300
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3388 25676 3444 25732
rect 9212 57708 9268 57764
rect 10892 70924 10948 70980
rect 7532 49532 7588 49588
rect 8428 46732 8484 46788
rect 10892 43372 10948 43428
rect 12908 66108 12964 66164
rect 10556 42812 10612 42868
rect 8428 37884 8484 37940
rect 8764 39676 8820 39732
rect 8764 35084 8820 35140
rect 7532 27244 7588 27300
rect 5852 25676 5908 25732
rect 9660 27020 9716 27076
rect 3500 24610 3556 24612
rect 3500 24558 3502 24610
rect 3502 24558 3554 24610
rect 3554 24558 3556 24610
rect 3500 24556 3556 24558
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3500 23042 3556 23044
rect 3500 22990 3502 23042
rect 3502 22990 3554 23042
rect 3554 22990 3556 23042
rect 3500 22988 3556 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4396 22146 4452 22148
rect 4396 22094 4398 22146
rect 4398 22094 4450 22146
rect 4450 22094 4452 22146
rect 4396 22092 4452 22094
rect 3612 21308 3668 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5628 19740 5684 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 3500 16882 3556 16884
rect 3500 16830 3502 16882
rect 3502 16830 3554 16882
rect 3554 16830 3556 16882
rect 3500 16828 3556 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 3052 10444 3108 10500
rect 1932 10220 1988 10276
rect 1820 6860 1876 6916
rect 1932 5516 1988 5572
rect 812 4396 868 4452
rect 140 3612 196 3668
rect 1932 4450 1988 4452
rect 1932 4398 1934 4450
rect 1934 4398 1986 4450
rect 1986 4398 1988 4450
rect 1932 4396 1988 4398
rect 1820 4172 1876 4228
rect 3052 6412 3108 6468
rect 3052 5906 3108 5908
rect 3052 5854 3054 5906
rect 3054 5854 3106 5906
rect 3106 5854 3108 5906
rect 3052 5852 3108 5854
rect 2380 4396 2436 4452
rect 2044 3612 2100 3668
rect 2156 4172 2212 4228
rect 2044 3442 2100 3444
rect 2044 3390 2046 3442
rect 2046 3390 2098 3442
rect 2098 3390 2100 3442
rect 2044 3388 2100 3390
rect 2828 4284 2884 4340
rect 3500 10498 3556 10500
rect 3500 10446 3502 10498
rect 3502 10446 3554 10498
rect 3554 10446 3556 10498
rect 3500 10444 3556 10446
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 3612 6466 3668 6468
rect 3612 6414 3614 6466
rect 3614 6414 3666 6466
rect 3666 6414 3668 6466
rect 3612 6412 3668 6414
rect 3500 5906 3556 5908
rect 3500 5854 3502 5906
rect 3502 5854 3554 5906
rect 3554 5854 3556 5906
rect 3500 5852 3556 5854
rect 3836 5740 3892 5796
rect 3164 4284 3220 4340
rect 3388 4396 3444 4452
rect 3724 3500 3780 3556
rect 2828 3388 2884 3444
rect 3500 3388 3556 3444
rect 5180 5794 5236 5796
rect 5180 5742 5182 5794
rect 5182 5742 5234 5794
rect 5234 5742 5236 5794
rect 5180 5740 5236 5742
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4956 5180 5012 5236
rect 4844 5122 4900 5124
rect 4844 5070 4846 5122
rect 4846 5070 4898 5122
rect 4898 5070 4900 5122
rect 4844 5068 4900 5070
rect 6076 5234 6132 5236
rect 6076 5182 6078 5234
rect 6078 5182 6130 5234
rect 6130 5182 6132 5234
rect 6076 5180 6132 5182
rect 5628 5068 5684 5124
rect 6524 5068 6580 5124
rect 3948 4226 4004 4228
rect 3948 4174 3950 4226
rect 3950 4174 4002 4226
rect 4002 4174 4004 4226
rect 3948 4172 4004 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4956 3666 5012 3668
rect 4956 3614 4958 3666
rect 4958 3614 5010 3666
rect 5010 3614 5012 3666
rect 4956 3612 5012 3614
rect 3500 2156 3556 2212
rect 6412 3388 6468 3444
rect 8204 4172 8260 4228
rect 8764 4226 8820 4228
rect 8764 4174 8766 4226
rect 8766 4174 8818 4226
rect 8818 4174 8820 4226
rect 8764 4172 8820 4174
rect 12348 31164 12404 31220
rect 12348 22988 12404 23044
rect 11228 4508 11284 4564
rect 11900 4562 11956 4564
rect 11900 4510 11902 4562
rect 11902 4510 11954 4562
rect 11954 4510 11956 4562
rect 11900 4508 11956 4510
rect 11228 4338 11284 4340
rect 11228 4286 11230 4338
rect 11230 4286 11282 4338
rect 11282 4286 11284 4338
rect 11228 4284 11284 4286
rect 11452 3612 11508 3668
rect 8876 3388 8932 3444
rect 9772 3442 9828 3444
rect 9772 3390 9774 3442
rect 9774 3390 9826 3442
rect 9826 3390 9828 3442
rect 9772 3388 9828 3390
rect 15932 97692 15988 97748
rect 17388 116450 17444 116452
rect 17388 116398 17390 116450
rect 17390 116398 17442 116450
rect 17442 116398 17444 116450
rect 17388 116396 17444 116398
rect 20972 116508 21028 116564
rect 19836 116058 19892 116060
rect 19836 116006 19838 116058
rect 19838 116006 19890 116058
rect 19890 116006 19892 116058
rect 19836 116004 19892 116006
rect 19940 116058 19996 116060
rect 19940 116006 19942 116058
rect 19942 116006 19994 116058
rect 19994 116006 19996 116058
rect 19940 116004 19996 116006
rect 20044 116058 20100 116060
rect 20044 116006 20046 116058
rect 20046 116006 20098 116058
rect 20098 116006 20100 116058
rect 20044 116004 20100 116006
rect 19836 114490 19892 114492
rect 19836 114438 19838 114490
rect 19838 114438 19890 114490
rect 19890 114438 19892 114490
rect 19836 114436 19892 114438
rect 19940 114490 19996 114492
rect 19940 114438 19942 114490
rect 19942 114438 19994 114490
rect 19994 114438 19996 114490
rect 19940 114436 19996 114438
rect 20044 114490 20100 114492
rect 20044 114438 20046 114490
rect 20046 114438 20098 114490
rect 20098 114438 20100 114490
rect 20044 114436 20100 114438
rect 19836 112922 19892 112924
rect 19836 112870 19838 112922
rect 19838 112870 19890 112922
rect 19890 112870 19892 112922
rect 19836 112868 19892 112870
rect 19940 112922 19996 112924
rect 19940 112870 19942 112922
rect 19942 112870 19994 112922
rect 19994 112870 19996 112922
rect 19940 112868 19996 112870
rect 20044 112922 20100 112924
rect 20044 112870 20046 112922
rect 20046 112870 20098 112922
rect 20098 112870 20100 112922
rect 20044 112868 20100 112870
rect 19836 111354 19892 111356
rect 19836 111302 19838 111354
rect 19838 111302 19890 111354
rect 19890 111302 19892 111354
rect 19836 111300 19892 111302
rect 19940 111354 19996 111356
rect 19940 111302 19942 111354
rect 19942 111302 19994 111354
rect 19994 111302 19996 111354
rect 19940 111300 19996 111302
rect 20044 111354 20100 111356
rect 20044 111302 20046 111354
rect 20046 111302 20098 111354
rect 20098 111302 20100 111354
rect 20044 111300 20100 111302
rect 19836 109786 19892 109788
rect 19836 109734 19838 109786
rect 19838 109734 19890 109786
rect 19890 109734 19892 109786
rect 19836 109732 19892 109734
rect 19940 109786 19996 109788
rect 19940 109734 19942 109786
rect 19942 109734 19994 109786
rect 19994 109734 19996 109786
rect 19940 109732 19996 109734
rect 20044 109786 20100 109788
rect 20044 109734 20046 109786
rect 20046 109734 20098 109786
rect 20098 109734 20100 109786
rect 20044 109732 20100 109734
rect 19836 108218 19892 108220
rect 19836 108166 19838 108218
rect 19838 108166 19890 108218
rect 19890 108166 19892 108218
rect 19836 108164 19892 108166
rect 19940 108218 19996 108220
rect 19940 108166 19942 108218
rect 19942 108166 19994 108218
rect 19994 108166 19996 108218
rect 19940 108164 19996 108166
rect 20044 108218 20100 108220
rect 20044 108166 20046 108218
rect 20046 108166 20098 108218
rect 20098 108166 20100 108218
rect 20044 108164 20100 108166
rect 19836 106650 19892 106652
rect 19836 106598 19838 106650
rect 19838 106598 19890 106650
rect 19890 106598 19892 106650
rect 19836 106596 19892 106598
rect 19940 106650 19996 106652
rect 19940 106598 19942 106650
rect 19942 106598 19994 106650
rect 19994 106598 19996 106650
rect 19940 106596 19996 106598
rect 20044 106650 20100 106652
rect 20044 106598 20046 106650
rect 20046 106598 20098 106650
rect 20098 106598 20100 106650
rect 20044 106596 20100 106598
rect 19836 105082 19892 105084
rect 19836 105030 19838 105082
rect 19838 105030 19890 105082
rect 19890 105030 19892 105082
rect 19836 105028 19892 105030
rect 19940 105082 19996 105084
rect 19940 105030 19942 105082
rect 19942 105030 19994 105082
rect 19994 105030 19996 105082
rect 19940 105028 19996 105030
rect 20044 105082 20100 105084
rect 20044 105030 20046 105082
rect 20046 105030 20098 105082
rect 20098 105030 20100 105082
rect 20044 105028 20100 105030
rect 19836 103514 19892 103516
rect 19836 103462 19838 103514
rect 19838 103462 19890 103514
rect 19890 103462 19892 103514
rect 19836 103460 19892 103462
rect 19940 103514 19996 103516
rect 19940 103462 19942 103514
rect 19942 103462 19994 103514
rect 19994 103462 19996 103514
rect 19940 103460 19996 103462
rect 20044 103514 20100 103516
rect 20044 103462 20046 103514
rect 20046 103462 20098 103514
rect 20098 103462 20100 103514
rect 20044 103460 20100 103462
rect 19836 101946 19892 101948
rect 19836 101894 19838 101946
rect 19838 101894 19890 101946
rect 19890 101894 19892 101946
rect 19836 101892 19892 101894
rect 19940 101946 19996 101948
rect 19940 101894 19942 101946
rect 19942 101894 19994 101946
rect 19994 101894 19996 101946
rect 19940 101892 19996 101894
rect 20044 101946 20100 101948
rect 20044 101894 20046 101946
rect 20046 101894 20098 101946
rect 20098 101894 20100 101946
rect 20044 101892 20100 101894
rect 19836 100378 19892 100380
rect 19836 100326 19838 100378
rect 19838 100326 19890 100378
rect 19890 100326 19892 100378
rect 19836 100324 19892 100326
rect 19940 100378 19996 100380
rect 19940 100326 19942 100378
rect 19942 100326 19994 100378
rect 19994 100326 19996 100378
rect 19940 100324 19996 100326
rect 20044 100378 20100 100380
rect 20044 100326 20046 100378
rect 20046 100326 20098 100378
rect 20098 100326 20100 100378
rect 20044 100324 20100 100326
rect 19836 98810 19892 98812
rect 19836 98758 19838 98810
rect 19838 98758 19890 98810
rect 19890 98758 19892 98810
rect 19836 98756 19892 98758
rect 19940 98810 19996 98812
rect 19940 98758 19942 98810
rect 19942 98758 19994 98810
rect 19994 98758 19996 98810
rect 19940 98756 19996 98758
rect 20044 98810 20100 98812
rect 20044 98758 20046 98810
rect 20046 98758 20098 98810
rect 20098 98758 20100 98810
rect 20044 98756 20100 98758
rect 19836 97242 19892 97244
rect 19836 97190 19838 97242
rect 19838 97190 19890 97242
rect 19890 97190 19892 97242
rect 19836 97188 19892 97190
rect 19940 97242 19996 97244
rect 19940 97190 19942 97242
rect 19942 97190 19994 97242
rect 19994 97190 19996 97242
rect 19940 97188 19996 97190
rect 20044 97242 20100 97244
rect 20044 97190 20046 97242
rect 20046 97190 20098 97242
rect 20098 97190 20100 97242
rect 20044 97188 20100 97190
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 16828 69916 16884 69972
rect 17612 69692 17668 69748
rect 15932 68012 15988 68068
rect 16156 68348 16212 68404
rect 14252 64652 14308 64708
rect 14252 48300 14308 48356
rect 13580 16828 13636 16884
rect 13580 15148 13636 15204
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 23548 116396 23604 116452
rect 22764 115890 22820 115892
rect 22764 115838 22766 115890
rect 22766 115838 22818 115890
rect 22818 115838 22820 115890
rect 22764 115836 22820 115838
rect 24332 116508 24388 116564
rect 26012 116562 26068 116564
rect 26012 116510 26014 116562
rect 26014 116510 26066 116562
rect 26066 116510 26068 116562
rect 26012 116508 26068 116510
rect 25340 116450 25396 116452
rect 25340 116398 25342 116450
rect 25342 116398 25394 116450
rect 25394 116398 25396 116450
rect 25340 116396 25396 116398
rect 24108 115890 24164 115892
rect 24108 115838 24110 115890
rect 24110 115838 24162 115890
rect 24162 115838 24164 115890
rect 24108 115836 24164 115838
rect 31500 116284 31556 116340
rect 23324 115666 23380 115668
rect 23324 115614 23326 115666
rect 23326 115614 23378 115666
rect 23378 115614 23380 115666
rect 23324 115612 23380 115614
rect 23324 114604 23380 114660
rect 23772 114658 23828 114660
rect 23772 114606 23774 114658
rect 23774 114606 23826 114658
rect 23826 114606 23828 114658
rect 23772 114604 23828 114606
rect 24668 114604 24724 114660
rect 29372 111804 29428 111860
rect 20972 63308 21028 63364
rect 22652 102396 22708 102452
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 22652 62300 22708 62356
rect 24332 88284 24388 88340
rect 24332 61292 24388 61348
rect 26012 76188 26068 76244
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 20972 59948 21028 60004
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 17612 56812 17668 56868
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 16156 47628 16212 47684
rect 17612 51212 17668 51268
rect 15932 42476 15988 42532
rect 15932 30156 15988 30212
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 17612 24556 17668 24612
rect 17836 23884 17892 23940
rect 14252 4396 14308 4452
rect 15372 9212 15428 9268
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 17836 5852 17892 5908
rect 19628 12684 19684 12740
rect 12908 3724 12964 3780
rect 12236 3666 12292 3668
rect 12236 3614 12238 3666
rect 12238 3614 12290 3666
rect 12290 3614 12292 3666
rect 12236 3612 12292 3614
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 26012 59276 26068 59332
rect 26012 57372 26068 57428
rect 22652 56700 22708 56756
rect 22652 41244 22708 41300
rect 24332 55020 24388 55076
rect 20972 5068 21028 5124
rect 22652 39788 22708 39844
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 16492 3666 16548 3668
rect 16492 3614 16494 3666
rect 16494 3614 16546 3666
rect 16546 3614 16548 3666
rect 16492 3612 16548 3614
rect 19628 3836 19684 3892
rect 20636 3724 20692 3780
rect 20972 3388 21028 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21532 3836 21588 3892
rect 33068 116338 33124 116340
rect 33068 116286 33070 116338
rect 33070 116286 33122 116338
rect 33122 116286 33124 116338
rect 33068 116284 33124 116286
rect 32844 115500 32900 115556
rect 33628 115554 33684 115556
rect 33628 115502 33630 115554
rect 33630 115502 33682 115554
rect 33682 115502 33684 115554
rect 33628 115500 33684 115502
rect 35196 116842 35252 116844
rect 35196 116790 35198 116842
rect 35198 116790 35250 116842
rect 35250 116790 35252 116842
rect 35196 116788 35252 116790
rect 35300 116842 35356 116844
rect 35300 116790 35302 116842
rect 35302 116790 35354 116842
rect 35354 116790 35356 116842
rect 35300 116788 35356 116790
rect 35404 116842 35460 116844
rect 35404 116790 35406 116842
rect 35406 116790 35458 116842
rect 35458 116790 35460 116842
rect 35404 116788 35460 116790
rect 35532 116508 35588 116564
rect 36316 115948 36372 116004
rect 37436 116562 37492 116564
rect 37436 116510 37438 116562
rect 37438 116510 37490 116562
rect 37490 116510 37492 116562
rect 37436 116508 37492 116510
rect 35196 115274 35252 115276
rect 35196 115222 35198 115274
rect 35198 115222 35250 115274
rect 35250 115222 35252 115274
rect 35196 115220 35252 115222
rect 35300 115274 35356 115276
rect 35300 115222 35302 115274
rect 35302 115222 35354 115274
rect 35354 115222 35356 115274
rect 35300 115220 35356 115222
rect 35404 115274 35460 115276
rect 35404 115222 35406 115274
rect 35406 115222 35458 115274
rect 35458 115222 35460 115274
rect 35404 115220 35460 115222
rect 33964 114604 34020 114660
rect 32172 101724 32228 101780
rect 32732 104524 32788 104580
rect 32732 66444 32788 66500
rect 32172 66332 32228 66388
rect 32172 59612 32228 59668
rect 33516 59052 33572 59108
rect 33516 55916 33572 55972
rect 30380 53452 30436 53508
rect 33516 54348 33572 54404
rect 29372 51548 29428 51604
rect 31052 52108 31108 52164
rect 27020 48860 27076 48916
rect 26012 22092 26068 22148
rect 26124 23660 26180 23716
rect 26124 10444 26180 10500
rect 24332 3612 24388 3668
rect 21196 3388 21252 3444
rect 21532 3442 21588 3444
rect 21532 3390 21534 3442
rect 21534 3390 21586 3442
rect 21586 3390 21588 3442
rect 21532 3388 21588 3390
rect 24668 3442 24724 3444
rect 24668 3390 24670 3442
rect 24670 3390 24722 3442
rect 24722 3390 24724 3442
rect 24668 3388 24724 3390
rect 26348 5122 26404 5124
rect 26348 5070 26350 5122
rect 26350 5070 26402 5122
rect 26402 5070 26404 5122
rect 26348 5068 26404 5070
rect 26908 5122 26964 5124
rect 26908 5070 26910 5122
rect 26910 5070 26962 5122
rect 26962 5070 26964 5122
rect 26908 5068 26964 5070
rect 25452 3442 25508 3444
rect 25452 3390 25454 3442
rect 25454 3390 25506 3442
rect 25506 3390 25508 3442
rect 25452 3388 25508 3390
rect 29372 44828 29428 44884
rect 29372 12684 29428 12740
rect 29484 26908 29540 26964
rect 29484 6412 29540 6468
rect 28140 5180 28196 5236
rect 34860 114604 34916 114660
rect 35532 114658 35588 114660
rect 35532 114606 35534 114658
rect 35534 114606 35586 114658
rect 35586 114606 35588 114658
rect 35532 114604 35588 114606
rect 35196 113706 35252 113708
rect 35196 113654 35198 113706
rect 35198 113654 35250 113706
rect 35250 113654 35252 113706
rect 35196 113652 35252 113654
rect 35300 113706 35356 113708
rect 35300 113654 35302 113706
rect 35302 113654 35354 113706
rect 35354 113654 35356 113706
rect 35300 113652 35356 113654
rect 35404 113706 35460 113708
rect 35404 113654 35406 113706
rect 35406 113654 35458 113706
rect 35458 113654 35460 113706
rect 35404 113652 35460 113654
rect 35196 112138 35252 112140
rect 35196 112086 35198 112138
rect 35198 112086 35250 112138
rect 35250 112086 35252 112138
rect 35196 112084 35252 112086
rect 35300 112138 35356 112140
rect 35300 112086 35302 112138
rect 35302 112086 35354 112138
rect 35354 112086 35356 112138
rect 35300 112084 35356 112086
rect 35404 112138 35460 112140
rect 35404 112086 35406 112138
rect 35406 112086 35458 112138
rect 35458 112086 35460 112138
rect 35404 112084 35460 112086
rect 35196 110570 35252 110572
rect 35196 110518 35198 110570
rect 35198 110518 35250 110570
rect 35250 110518 35252 110570
rect 35196 110516 35252 110518
rect 35300 110570 35356 110572
rect 35300 110518 35302 110570
rect 35302 110518 35354 110570
rect 35354 110518 35356 110570
rect 35300 110516 35356 110518
rect 35404 110570 35460 110572
rect 35404 110518 35406 110570
rect 35406 110518 35458 110570
rect 35458 110518 35460 110570
rect 35404 110516 35460 110518
rect 35196 109002 35252 109004
rect 35196 108950 35198 109002
rect 35198 108950 35250 109002
rect 35250 108950 35252 109002
rect 35196 108948 35252 108950
rect 35300 109002 35356 109004
rect 35300 108950 35302 109002
rect 35302 108950 35354 109002
rect 35354 108950 35356 109002
rect 35300 108948 35356 108950
rect 35404 109002 35460 109004
rect 35404 108950 35406 109002
rect 35406 108950 35458 109002
rect 35458 108950 35460 109002
rect 35404 108948 35460 108950
rect 35196 107434 35252 107436
rect 35196 107382 35198 107434
rect 35198 107382 35250 107434
rect 35250 107382 35252 107434
rect 35196 107380 35252 107382
rect 35300 107434 35356 107436
rect 35300 107382 35302 107434
rect 35302 107382 35354 107434
rect 35354 107382 35356 107434
rect 35300 107380 35356 107382
rect 35404 107434 35460 107436
rect 35404 107382 35406 107434
rect 35406 107382 35458 107434
rect 35458 107382 35460 107434
rect 35404 107380 35460 107382
rect 35196 105866 35252 105868
rect 35196 105814 35198 105866
rect 35198 105814 35250 105866
rect 35250 105814 35252 105866
rect 35196 105812 35252 105814
rect 35300 105866 35356 105868
rect 35300 105814 35302 105866
rect 35302 105814 35354 105866
rect 35354 105814 35356 105866
rect 35300 105812 35356 105814
rect 35404 105866 35460 105868
rect 35404 105814 35406 105866
rect 35406 105814 35458 105866
rect 35458 105814 35460 105866
rect 35404 105812 35460 105814
rect 35196 104298 35252 104300
rect 35196 104246 35198 104298
rect 35198 104246 35250 104298
rect 35250 104246 35252 104298
rect 35196 104244 35252 104246
rect 35300 104298 35356 104300
rect 35300 104246 35302 104298
rect 35302 104246 35354 104298
rect 35354 104246 35356 104298
rect 35300 104244 35356 104246
rect 35404 104298 35460 104300
rect 35404 104246 35406 104298
rect 35406 104246 35458 104298
rect 35458 104246 35460 104298
rect 35404 104244 35460 104246
rect 35196 102730 35252 102732
rect 35196 102678 35198 102730
rect 35198 102678 35250 102730
rect 35250 102678 35252 102730
rect 35196 102676 35252 102678
rect 35300 102730 35356 102732
rect 35300 102678 35302 102730
rect 35302 102678 35354 102730
rect 35354 102678 35356 102730
rect 35300 102676 35356 102678
rect 35404 102730 35460 102732
rect 35404 102678 35406 102730
rect 35406 102678 35458 102730
rect 35458 102678 35460 102730
rect 35404 102676 35460 102678
rect 35196 101162 35252 101164
rect 35196 101110 35198 101162
rect 35198 101110 35250 101162
rect 35250 101110 35252 101162
rect 35196 101108 35252 101110
rect 35300 101162 35356 101164
rect 35300 101110 35302 101162
rect 35302 101110 35354 101162
rect 35354 101110 35356 101162
rect 35300 101108 35356 101110
rect 35404 101162 35460 101164
rect 35404 101110 35406 101162
rect 35406 101110 35458 101162
rect 35458 101110 35460 101162
rect 35404 101108 35460 101110
rect 35196 99594 35252 99596
rect 35196 99542 35198 99594
rect 35198 99542 35250 99594
rect 35250 99542 35252 99594
rect 35196 99540 35252 99542
rect 35300 99594 35356 99596
rect 35300 99542 35302 99594
rect 35302 99542 35354 99594
rect 35354 99542 35356 99594
rect 35300 99540 35356 99542
rect 35404 99594 35460 99596
rect 35404 99542 35406 99594
rect 35406 99542 35458 99594
rect 35458 99542 35460 99594
rect 35404 99540 35460 99542
rect 35196 98026 35252 98028
rect 35196 97974 35198 98026
rect 35198 97974 35250 98026
rect 35250 97974 35252 98026
rect 35196 97972 35252 97974
rect 35300 98026 35356 98028
rect 35300 97974 35302 98026
rect 35302 97974 35354 98026
rect 35354 97974 35356 98026
rect 35300 97972 35356 97974
rect 35404 98026 35460 98028
rect 35404 97974 35406 98026
rect 35406 97974 35458 98026
rect 35458 97974 35460 98026
rect 35404 97972 35460 97974
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 37772 115500 37828 115556
rect 36652 66332 36708 66388
rect 36876 69916 36932 69972
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 36876 65100 36932 65156
rect 35404 65044 35460 65046
rect 36316 64652 36372 64708
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 38668 115554 38724 115556
rect 38668 115502 38670 115554
rect 38670 115502 38722 115554
rect 38722 115502 38724 115554
rect 38668 115500 38724 115502
rect 43148 116284 43204 116340
rect 43484 116396 43540 116452
rect 42140 115948 42196 116004
rect 41132 115500 41188 115556
rect 37884 99820 37940 99876
rect 38556 99426 38612 99428
rect 38556 99374 38558 99426
rect 38558 99374 38610 99426
rect 38610 99374 38612 99426
rect 38556 99372 38612 99374
rect 39452 99372 39508 99428
rect 39564 101724 39620 101780
rect 38892 99202 38948 99204
rect 38892 99150 38894 99202
rect 38894 99150 38946 99202
rect 38946 99150 38948 99202
rect 38892 99148 38948 99150
rect 37772 63980 37828 64036
rect 36316 57596 36372 57652
rect 37772 60172 37828 60228
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 36204 56364 36260 56420
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 33516 52108 33572 52164
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34412 51100 34468 51156
rect 34636 51100 34692 51156
rect 32732 47516 32788 47572
rect 32732 41132 32788 41188
rect 32172 40348 32228 40404
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36092 40236 36148 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34636 31164 34692 31220
rect 34412 31052 34468 31108
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34524 21420 34580 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34524 5180 34580 5236
rect 37548 41692 37604 41748
rect 42140 113372 42196 113428
rect 41692 99148 41748 99204
rect 40012 55410 40068 55412
rect 40012 55358 40014 55410
rect 40014 55358 40066 55410
rect 40066 55358 40068 55410
rect 40012 55356 40068 55358
rect 40908 55356 40964 55412
rect 40796 55298 40852 55300
rect 40796 55246 40798 55298
rect 40798 55246 40850 55298
rect 40850 55246 40852 55298
rect 40796 55244 40852 55246
rect 39676 55074 39732 55076
rect 39676 55022 39678 55074
rect 39678 55022 39730 55074
rect 39730 55022 39732 55074
rect 39676 55020 39732 55022
rect 40684 55074 40740 55076
rect 40684 55022 40686 55074
rect 40686 55022 40738 55074
rect 40738 55022 40740 55074
rect 40684 55020 40740 55022
rect 40908 54572 40964 54628
rect 40348 54402 40404 54404
rect 40348 54350 40350 54402
rect 40350 54350 40402 54402
rect 40402 54350 40404 54402
rect 40348 54348 40404 54350
rect 39564 50316 39620 50372
rect 37772 40348 37828 40404
rect 39116 48748 39172 48804
rect 37548 36540 37604 36596
rect 36204 32396 36260 32452
rect 37772 33404 37828 33460
rect 37772 9212 37828 9268
rect 36092 5068 36148 5124
rect 36540 4060 36596 4116
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34412 3724 34468 3780
rect 41692 55804 41748 55860
rect 42252 55020 42308 55076
rect 43372 55020 43428 55076
rect 41580 54626 41636 54628
rect 41580 54574 41582 54626
rect 41582 54574 41634 54626
rect 41634 54574 41636 54626
rect 41580 54572 41636 54574
rect 41804 54348 41860 54404
rect 42476 53788 42532 53844
rect 43372 53788 43428 53844
rect 42028 51996 42084 52052
rect 43148 51996 43204 52052
rect 43372 51996 43428 52052
rect 43596 116060 43652 116116
rect 44044 116338 44100 116340
rect 44044 116286 44046 116338
rect 44046 116286 44098 116338
rect 44098 116286 44100 116338
rect 44044 116284 44100 116286
rect 46956 116338 47012 116340
rect 46956 116286 46958 116338
rect 46958 116286 47010 116338
rect 47010 116286 47012 116338
rect 46956 116284 47012 116286
rect 47628 116284 47684 116340
rect 48748 116338 48804 116340
rect 48748 116286 48750 116338
rect 48750 116286 48802 116338
rect 48802 116286 48804 116338
rect 48748 116284 48804 116286
rect 51212 116396 51268 116452
rect 48076 116172 48132 116228
rect 48524 116060 48580 116116
rect 46508 115724 46564 115780
rect 47964 115724 48020 115780
rect 43596 114940 43652 114996
rect 45388 114994 45444 114996
rect 45388 114942 45390 114994
rect 45390 114942 45442 114994
rect 45442 114942 45444 114994
rect 45388 114940 45444 114942
rect 46396 114940 46452 114996
rect 45276 105756 45332 105812
rect 44828 102956 44884 103012
rect 45164 102956 45220 103012
rect 44604 66444 44660 66500
rect 44716 64540 44772 64596
rect 44492 58156 44548 58212
rect 45612 103010 45668 103012
rect 45612 102958 45614 103010
rect 45614 102958 45666 103010
rect 45666 102958 45668 103010
rect 45612 102956 45668 102958
rect 45948 102956 46004 103012
rect 46956 114994 47012 114996
rect 46956 114942 46958 114994
rect 46958 114942 47010 114994
rect 47010 114942 47012 114994
rect 46956 114940 47012 114942
rect 46508 105756 46564 105812
rect 48300 93548 48356 93604
rect 46060 68460 46116 68516
rect 46844 68514 46900 68516
rect 46844 68462 46846 68514
rect 46846 68462 46898 68514
rect 46898 68462 46900 68514
rect 46844 68460 46900 68462
rect 45612 63868 45668 63924
rect 46396 66668 46452 66724
rect 45836 65548 45892 65604
rect 45948 64706 46004 64708
rect 45948 64654 45950 64706
rect 45950 64654 46002 64706
rect 46002 64654 46004 64706
rect 45948 64652 46004 64654
rect 45836 63980 45892 64036
rect 45724 63532 45780 63588
rect 46732 65602 46788 65604
rect 46732 65550 46734 65602
rect 46734 65550 46786 65602
rect 46786 65550 46788 65602
rect 46732 65548 46788 65550
rect 46732 64876 46788 64932
rect 48412 67058 48468 67060
rect 48412 67006 48414 67058
rect 48414 67006 48466 67058
rect 48466 67006 48468 67058
rect 48412 67004 48468 67006
rect 47964 66892 48020 66948
rect 47292 66386 47348 66388
rect 47292 66334 47294 66386
rect 47294 66334 47346 66386
rect 47346 66334 47348 66386
rect 47292 66332 47348 66334
rect 47516 65490 47572 65492
rect 47516 65438 47518 65490
rect 47518 65438 47570 65490
rect 47570 65438 47572 65490
rect 47516 65436 47572 65438
rect 46844 64764 46900 64820
rect 47628 64876 47684 64932
rect 47180 64652 47236 64708
rect 46508 64594 46564 64596
rect 46508 64542 46510 64594
rect 46510 64542 46562 64594
rect 46562 64542 46564 64594
rect 46508 64540 46564 64542
rect 46844 64540 46900 64596
rect 46060 60786 46116 60788
rect 46060 60734 46062 60786
rect 46062 60734 46114 60786
rect 46114 60734 46116 60786
rect 46060 60732 46116 60734
rect 45276 60060 45332 60116
rect 44604 57260 44660 57316
rect 46620 59836 46676 59892
rect 44492 56252 44548 56308
rect 44940 56588 44996 56644
rect 46172 56140 46228 56196
rect 44940 54684 44996 54740
rect 45612 55916 45668 55972
rect 45388 53618 45444 53620
rect 45388 53566 45390 53618
rect 45390 53566 45442 53618
rect 45442 53566 45444 53618
rect 45388 53564 45444 53566
rect 45052 51490 45108 51492
rect 45052 51438 45054 51490
rect 45054 51438 45106 51490
rect 45106 51438 45108 51490
rect 45052 51436 45108 51438
rect 45388 51436 45444 51492
rect 45500 51100 45556 51156
rect 45724 54738 45780 54740
rect 45724 54686 45726 54738
rect 45726 54686 45778 54738
rect 45778 54686 45780 54738
rect 45724 54684 45780 54686
rect 45724 54460 45780 54516
rect 46172 54626 46228 54628
rect 46172 54574 46174 54626
rect 46174 54574 46226 54626
rect 46226 54574 46228 54626
rect 46172 54572 46228 54574
rect 46508 54796 46564 54852
rect 46508 54572 46564 54628
rect 45948 53730 46004 53732
rect 45948 53678 45950 53730
rect 45950 53678 46002 53730
rect 46002 53678 46004 53730
rect 45948 53676 46004 53678
rect 46060 52274 46116 52276
rect 46060 52222 46062 52274
rect 46062 52222 46114 52274
rect 46114 52222 46116 52274
rect 46060 52220 46116 52222
rect 45836 51324 45892 51380
rect 46060 50876 46116 50932
rect 45836 50540 45892 50596
rect 47068 60732 47124 60788
rect 47068 56194 47124 56196
rect 47068 56142 47070 56194
rect 47070 56142 47122 56194
rect 47122 56142 47124 56194
rect 47068 56140 47124 56142
rect 46956 56028 47012 56084
rect 45500 49810 45556 49812
rect 45500 49758 45502 49810
rect 45502 49758 45554 49810
rect 45554 49758 45556 49810
rect 45500 49756 45556 49758
rect 45276 49644 45332 49700
rect 43484 48412 43540 48468
rect 45724 48972 45780 49028
rect 45724 48802 45780 48804
rect 45724 48750 45726 48802
rect 45726 48750 45778 48802
rect 45778 48750 45780 48802
rect 45724 48748 45780 48750
rect 45724 48300 45780 48356
rect 41244 47740 41300 47796
rect 45500 47570 45556 47572
rect 45500 47518 45502 47570
rect 45502 47518 45554 47570
rect 45554 47518 45556 47570
rect 45500 47516 45556 47518
rect 42924 46172 42980 46228
rect 42140 45218 42196 45220
rect 42140 45166 42142 45218
rect 42142 45166 42194 45218
rect 42194 45166 42196 45218
rect 42140 45164 42196 45166
rect 43596 45500 43652 45556
rect 41916 45052 41972 45108
rect 41132 43148 41188 43204
rect 39452 21308 39508 21364
rect 39788 20860 39844 20916
rect 40236 20914 40292 20916
rect 40236 20862 40238 20914
rect 40238 20862 40290 20914
rect 40290 20862 40292 20914
rect 40236 20860 40292 20862
rect 41916 42812 41972 42868
rect 41132 20860 41188 20916
rect 43148 40572 43204 40628
rect 41580 5180 41636 5236
rect 42028 4508 42084 4564
rect 42364 5010 42420 5012
rect 42364 4958 42366 5010
rect 42366 4958 42418 5010
rect 42418 4958 42420 5010
rect 42364 4956 42420 4958
rect 42364 4508 42420 4564
rect 45612 45052 45668 45108
rect 44940 41804 44996 41860
rect 45836 40290 45892 40292
rect 45836 40238 45838 40290
rect 45838 40238 45890 40290
rect 45890 40238 45892 40290
rect 45836 40236 45892 40238
rect 46396 51324 46452 51380
rect 46396 50428 46452 50484
rect 46396 50316 46452 50372
rect 47068 54402 47124 54404
rect 47068 54350 47070 54402
rect 47070 54350 47122 54402
rect 47122 54350 47124 54402
rect 47068 54348 47124 54350
rect 46844 53900 46900 53956
rect 47964 64876 48020 64932
rect 47852 64594 47908 64596
rect 47852 64542 47854 64594
rect 47854 64542 47906 64594
rect 47906 64542 47908 64594
rect 47852 64540 47908 64542
rect 48188 64428 48244 64484
rect 48412 63756 48468 63812
rect 48188 63644 48244 63700
rect 48076 62412 48132 62468
rect 47740 62076 47796 62132
rect 47404 59890 47460 59892
rect 47404 59838 47406 59890
rect 47406 59838 47458 59890
rect 47458 59838 47460 59890
rect 47404 59836 47460 59838
rect 47964 60114 48020 60116
rect 47964 60062 47966 60114
rect 47966 60062 48018 60114
rect 48018 60062 48020 60114
rect 47964 60060 48020 60062
rect 47404 56866 47460 56868
rect 47404 56814 47406 56866
rect 47406 56814 47458 56866
rect 47458 56814 47460 56866
rect 47404 56812 47460 56814
rect 47852 56082 47908 56084
rect 47852 56030 47854 56082
rect 47854 56030 47906 56082
rect 47906 56030 47908 56082
rect 47852 56028 47908 56030
rect 47964 55692 48020 55748
rect 48300 62076 48356 62132
rect 50556 116058 50612 116060
rect 50556 116006 50558 116058
rect 50558 116006 50610 116058
rect 50610 116006 50612 116058
rect 50556 116004 50612 116006
rect 50660 116058 50716 116060
rect 50660 116006 50662 116058
rect 50662 116006 50714 116058
rect 50714 116006 50716 116058
rect 50660 116004 50716 116006
rect 50764 116058 50820 116060
rect 50764 116006 50766 116058
rect 50766 116006 50818 116058
rect 50818 116006 50820 116058
rect 50764 116004 50820 116006
rect 52108 116620 52164 116676
rect 53228 116508 53284 116564
rect 54012 116562 54068 116564
rect 54012 116510 54014 116562
rect 54014 116510 54066 116562
rect 54066 116510 54068 116562
rect 54012 116508 54068 116510
rect 52108 115948 52164 116004
rect 50556 114490 50612 114492
rect 50556 114438 50558 114490
rect 50558 114438 50610 114490
rect 50610 114438 50612 114490
rect 50556 114436 50612 114438
rect 50660 114490 50716 114492
rect 50660 114438 50662 114490
rect 50662 114438 50714 114490
rect 50714 114438 50716 114490
rect 50660 114436 50716 114438
rect 50764 114490 50820 114492
rect 50764 114438 50766 114490
rect 50766 114438 50818 114490
rect 50818 114438 50820 114490
rect 50764 114436 50820 114438
rect 50556 112922 50612 112924
rect 50556 112870 50558 112922
rect 50558 112870 50610 112922
rect 50610 112870 50612 112922
rect 50556 112868 50612 112870
rect 50660 112922 50716 112924
rect 50660 112870 50662 112922
rect 50662 112870 50714 112922
rect 50714 112870 50716 112922
rect 50660 112868 50716 112870
rect 50764 112922 50820 112924
rect 50764 112870 50766 112922
rect 50766 112870 50818 112922
rect 50818 112870 50820 112922
rect 50764 112868 50820 112870
rect 50556 111354 50612 111356
rect 50556 111302 50558 111354
rect 50558 111302 50610 111354
rect 50610 111302 50612 111354
rect 50556 111300 50612 111302
rect 50660 111354 50716 111356
rect 50660 111302 50662 111354
rect 50662 111302 50714 111354
rect 50714 111302 50716 111354
rect 50660 111300 50716 111302
rect 50764 111354 50820 111356
rect 50764 111302 50766 111354
rect 50766 111302 50818 111354
rect 50818 111302 50820 111354
rect 50764 111300 50820 111302
rect 50556 109786 50612 109788
rect 50556 109734 50558 109786
rect 50558 109734 50610 109786
rect 50610 109734 50612 109786
rect 50556 109732 50612 109734
rect 50660 109786 50716 109788
rect 50660 109734 50662 109786
rect 50662 109734 50714 109786
rect 50714 109734 50716 109786
rect 50660 109732 50716 109734
rect 50764 109786 50820 109788
rect 50764 109734 50766 109786
rect 50766 109734 50818 109786
rect 50818 109734 50820 109786
rect 50764 109732 50820 109734
rect 50556 108218 50612 108220
rect 50556 108166 50558 108218
rect 50558 108166 50610 108218
rect 50610 108166 50612 108218
rect 50556 108164 50612 108166
rect 50660 108218 50716 108220
rect 50660 108166 50662 108218
rect 50662 108166 50714 108218
rect 50714 108166 50716 108218
rect 50660 108164 50716 108166
rect 50764 108218 50820 108220
rect 50764 108166 50766 108218
rect 50766 108166 50818 108218
rect 50818 108166 50820 108218
rect 50764 108164 50820 108166
rect 50556 106650 50612 106652
rect 50556 106598 50558 106650
rect 50558 106598 50610 106650
rect 50610 106598 50612 106650
rect 50556 106596 50612 106598
rect 50660 106650 50716 106652
rect 50660 106598 50662 106650
rect 50662 106598 50714 106650
rect 50714 106598 50716 106650
rect 50660 106596 50716 106598
rect 50764 106650 50820 106652
rect 50764 106598 50766 106650
rect 50766 106598 50818 106650
rect 50818 106598 50820 106650
rect 50764 106596 50820 106598
rect 52444 105196 52500 105252
rect 50556 105082 50612 105084
rect 50556 105030 50558 105082
rect 50558 105030 50610 105082
rect 50610 105030 50612 105082
rect 50556 105028 50612 105030
rect 50660 105082 50716 105084
rect 50660 105030 50662 105082
rect 50662 105030 50714 105082
rect 50714 105030 50716 105082
rect 50660 105028 50716 105030
rect 50764 105082 50820 105084
rect 50764 105030 50766 105082
rect 50766 105030 50818 105082
rect 50818 105030 50820 105082
rect 50764 105028 50820 105030
rect 50556 103514 50612 103516
rect 50556 103462 50558 103514
rect 50558 103462 50610 103514
rect 50610 103462 50612 103514
rect 50556 103460 50612 103462
rect 50660 103514 50716 103516
rect 50660 103462 50662 103514
rect 50662 103462 50714 103514
rect 50714 103462 50716 103514
rect 50660 103460 50716 103462
rect 50764 103514 50820 103516
rect 50764 103462 50766 103514
rect 50766 103462 50818 103514
rect 50818 103462 50820 103514
rect 50764 103460 50820 103462
rect 50556 101946 50612 101948
rect 50556 101894 50558 101946
rect 50558 101894 50610 101946
rect 50610 101894 50612 101946
rect 50556 101892 50612 101894
rect 50660 101946 50716 101948
rect 50660 101894 50662 101946
rect 50662 101894 50714 101946
rect 50714 101894 50716 101946
rect 50660 101892 50716 101894
rect 50764 101946 50820 101948
rect 50764 101894 50766 101946
rect 50766 101894 50818 101946
rect 50818 101894 50820 101946
rect 50764 101892 50820 101894
rect 50556 100378 50612 100380
rect 50556 100326 50558 100378
rect 50558 100326 50610 100378
rect 50610 100326 50612 100378
rect 50556 100324 50612 100326
rect 50660 100378 50716 100380
rect 50660 100326 50662 100378
rect 50662 100326 50714 100378
rect 50714 100326 50716 100378
rect 50660 100324 50716 100326
rect 50764 100378 50820 100380
rect 50764 100326 50766 100378
rect 50766 100326 50818 100378
rect 50818 100326 50820 100378
rect 50764 100324 50820 100326
rect 50556 98810 50612 98812
rect 50556 98758 50558 98810
rect 50558 98758 50610 98810
rect 50610 98758 50612 98810
rect 50556 98756 50612 98758
rect 50660 98810 50716 98812
rect 50660 98758 50662 98810
rect 50662 98758 50714 98810
rect 50714 98758 50716 98810
rect 50660 98756 50716 98758
rect 50764 98810 50820 98812
rect 50764 98758 50766 98810
rect 50766 98758 50818 98810
rect 50818 98758 50820 98810
rect 50764 98756 50820 98758
rect 50556 97242 50612 97244
rect 50556 97190 50558 97242
rect 50558 97190 50610 97242
rect 50610 97190 50612 97242
rect 50556 97188 50612 97190
rect 50660 97242 50716 97244
rect 50660 97190 50662 97242
rect 50662 97190 50714 97242
rect 50714 97190 50716 97242
rect 50660 97188 50716 97190
rect 50764 97242 50820 97244
rect 50764 97190 50766 97242
rect 50766 97190 50818 97242
rect 50818 97190 50820 97242
rect 50764 97188 50820 97190
rect 50556 95674 50612 95676
rect 50556 95622 50558 95674
rect 50558 95622 50610 95674
rect 50610 95622 50612 95674
rect 50556 95620 50612 95622
rect 50660 95674 50716 95676
rect 50660 95622 50662 95674
rect 50662 95622 50714 95674
rect 50714 95622 50716 95674
rect 50660 95620 50716 95622
rect 50764 95674 50820 95676
rect 50764 95622 50766 95674
rect 50766 95622 50818 95674
rect 50818 95622 50820 95674
rect 50764 95620 50820 95622
rect 50556 94106 50612 94108
rect 50556 94054 50558 94106
rect 50558 94054 50610 94106
rect 50610 94054 50612 94106
rect 50556 94052 50612 94054
rect 50660 94106 50716 94108
rect 50660 94054 50662 94106
rect 50662 94054 50714 94106
rect 50714 94054 50716 94106
rect 50660 94052 50716 94054
rect 50764 94106 50820 94108
rect 50764 94054 50766 94106
rect 50766 94054 50818 94106
rect 50818 94054 50820 94106
rect 50764 94052 50820 94054
rect 48636 93548 48692 93604
rect 49420 93602 49476 93604
rect 49420 93550 49422 93602
rect 49422 93550 49474 93602
rect 49474 93550 49476 93602
rect 49420 93548 49476 93550
rect 50556 92538 50612 92540
rect 50556 92486 50558 92538
rect 50558 92486 50610 92538
rect 50610 92486 50612 92538
rect 50556 92484 50612 92486
rect 50660 92538 50716 92540
rect 50660 92486 50662 92538
rect 50662 92486 50714 92538
rect 50714 92486 50716 92538
rect 50660 92484 50716 92486
rect 50764 92538 50820 92540
rect 50764 92486 50766 92538
rect 50766 92486 50818 92538
rect 50818 92486 50820 92538
rect 50764 92484 50820 92486
rect 50556 90970 50612 90972
rect 50556 90918 50558 90970
rect 50558 90918 50610 90970
rect 50610 90918 50612 90970
rect 50556 90916 50612 90918
rect 50660 90970 50716 90972
rect 50660 90918 50662 90970
rect 50662 90918 50714 90970
rect 50714 90918 50716 90970
rect 50660 90916 50716 90918
rect 50764 90970 50820 90972
rect 50764 90918 50766 90970
rect 50766 90918 50818 90970
rect 50818 90918 50820 90970
rect 50764 90916 50820 90918
rect 50556 89402 50612 89404
rect 50556 89350 50558 89402
rect 50558 89350 50610 89402
rect 50610 89350 50612 89402
rect 50556 89348 50612 89350
rect 50660 89402 50716 89404
rect 50660 89350 50662 89402
rect 50662 89350 50714 89402
rect 50714 89350 50716 89402
rect 50660 89348 50716 89350
rect 50764 89402 50820 89404
rect 50764 89350 50766 89402
rect 50766 89350 50818 89402
rect 50818 89350 50820 89402
rect 50764 89348 50820 89350
rect 50556 87834 50612 87836
rect 50556 87782 50558 87834
rect 50558 87782 50610 87834
rect 50610 87782 50612 87834
rect 50556 87780 50612 87782
rect 50660 87834 50716 87836
rect 50660 87782 50662 87834
rect 50662 87782 50714 87834
rect 50714 87782 50716 87834
rect 50660 87780 50716 87782
rect 50764 87834 50820 87836
rect 50764 87782 50766 87834
rect 50766 87782 50818 87834
rect 50818 87782 50820 87834
rect 50764 87780 50820 87782
rect 50556 86266 50612 86268
rect 50556 86214 50558 86266
rect 50558 86214 50610 86266
rect 50610 86214 50612 86266
rect 50556 86212 50612 86214
rect 50660 86266 50716 86268
rect 50660 86214 50662 86266
rect 50662 86214 50714 86266
rect 50714 86214 50716 86266
rect 50660 86212 50716 86214
rect 50764 86266 50820 86268
rect 50764 86214 50766 86266
rect 50766 86214 50818 86266
rect 50818 86214 50820 86266
rect 50764 86212 50820 86214
rect 50556 84698 50612 84700
rect 50556 84646 50558 84698
rect 50558 84646 50610 84698
rect 50610 84646 50612 84698
rect 50556 84644 50612 84646
rect 50660 84698 50716 84700
rect 50660 84646 50662 84698
rect 50662 84646 50714 84698
rect 50714 84646 50716 84698
rect 50660 84644 50716 84646
rect 50764 84698 50820 84700
rect 50764 84646 50766 84698
rect 50766 84646 50818 84698
rect 50818 84646 50820 84698
rect 50764 84644 50820 84646
rect 50556 83130 50612 83132
rect 50556 83078 50558 83130
rect 50558 83078 50610 83130
rect 50610 83078 50612 83130
rect 50556 83076 50612 83078
rect 50660 83130 50716 83132
rect 50660 83078 50662 83130
rect 50662 83078 50714 83130
rect 50714 83078 50716 83130
rect 50660 83076 50716 83078
rect 50764 83130 50820 83132
rect 50764 83078 50766 83130
rect 50766 83078 50818 83130
rect 50818 83078 50820 83130
rect 50764 83076 50820 83078
rect 50556 81562 50612 81564
rect 50556 81510 50558 81562
rect 50558 81510 50610 81562
rect 50610 81510 50612 81562
rect 50556 81508 50612 81510
rect 50660 81562 50716 81564
rect 50660 81510 50662 81562
rect 50662 81510 50714 81562
rect 50714 81510 50716 81562
rect 50660 81508 50716 81510
rect 50764 81562 50820 81564
rect 50764 81510 50766 81562
rect 50766 81510 50818 81562
rect 50818 81510 50820 81562
rect 50764 81508 50820 81510
rect 50556 79994 50612 79996
rect 50556 79942 50558 79994
rect 50558 79942 50610 79994
rect 50610 79942 50612 79994
rect 50556 79940 50612 79942
rect 50660 79994 50716 79996
rect 50660 79942 50662 79994
rect 50662 79942 50714 79994
rect 50714 79942 50716 79994
rect 50660 79940 50716 79942
rect 50764 79994 50820 79996
rect 50764 79942 50766 79994
rect 50766 79942 50818 79994
rect 50818 79942 50820 79994
rect 50764 79940 50820 79942
rect 50556 78426 50612 78428
rect 50556 78374 50558 78426
rect 50558 78374 50610 78426
rect 50610 78374 50612 78426
rect 50556 78372 50612 78374
rect 50660 78426 50716 78428
rect 50660 78374 50662 78426
rect 50662 78374 50714 78426
rect 50714 78374 50716 78426
rect 50660 78372 50716 78374
rect 50764 78426 50820 78428
rect 50764 78374 50766 78426
rect 50766 78374 50818 78426
rect 50818 78374 50820 78426
rect 50764 78372 50820 78374
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 49532 67116 49588 67172
rect 49644 67058 49700 67060
rect 49644 67006 49646 67058
rect 49646 67006 49698 67058
rect 49698 67006 49700 67058
rect 49644 67004 49700 67006
rect 49532 66444 49588 66500
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 50540 67170 50596 67172
rect 50540 67118 50542 67170
rect 50542 67118 50594 67170
rect 50594 67118 50596 67170
rect 50540 67116 50596 67118
rect 51996 67004 52052 67060
rect 50764 66892 50820 66948
rect 48636 66332 48692 66388
rect 49420 66386 49476 66388
rect 49420 66334 49422 66386
rect 49422 66334 49474 66386
rect 49474 66334 49476 66386
rect 49420 66332 49476 66334
rect 48636 65436 48692 65492
rect 49532 65490 49588 65492
rect 49532 65438 49534 65490
rect 49534 65438 49586 65490
rect 49586 65438 49588 65490
rect 49532 65436 49588 65438
rect 48748 65212 48804 65268
rect 48748 64540 48804 64596
rect 48636 63922 48692 63924
rect 48636 63870 48638 63922
rect 48638 63870 48690 63922
rect 48690 63870 48692 63922
rect 48636 63868 48692 63870
rect 48636 63250 48692 63252
rect 48636 63198 48638 63250
rect 48638 63198 48690 63250
rect 48690 63198 48692 63250
rect 48636 63196 48692 63198
rect 48524 61964 48580 62020
rect 49644 64034 49700 64036
rect 49644 63982 49646 64034
rect 49646 63982 49698 64034
rect 49698 63982 49700 64034
rect 49644 63980 49700 63982
rect 49532 63810 49588 63812
rect 49532 63758 49534 63810
rect 49534 63758 49586 63810
rect 49586 63758 49588 63810
rect 49532 63756 49588 63758
rect 49196 62412 49252 62468
rect 49532 62466 49588 62468
rect 49532 62414 49534 62466
rect 49534 62414 49586 62466
rect 49586 62414 49588 62466
rect 49532 62412 49588 62414
rect 50764 66668 50820 66724
rect 51324 66668 51380 66724
rect 50652 66050 50708 66052
rect 50652 65998 50654 66050
rect 50654 65998 50706 66050
rect 50706 65998 50708 66050
rect 50652 65996 50708 65998
rect 51884 66108 51940 66164
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 49980 65490 50036 65492
rect 49980 65438 49982 65490
rect 49982 65438 50034 65490
rect 50034 65438 50036 65490
rect 49980 65436 50036 65438
rect 50652 64482 50708 64484
rect 50652 64430 50654 64482
rect 50654 64430 50706 64482
rect 50706 64430 50708 64482
rect 50652 64428 50708 64430
rect 51436 64428 51492 64484
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50428 63810 50484 63812
rect 50428 63758 50430 63810
rect 50430 63758 50482 63810
rect 50482 63758 50484 63810
rect 50428 63756 50484 63758
rect 50204 63644 50260 63700
rect 49868 62860 49924 62916
rect 50764 63196 50820 63252
rect 50316 62972 50372 63028
rect 50764 63026 50820 63028
rect 50764 62974 50766 63026
rect 50766 62974 50818 63026
rect 50818 62974 50820 63026
rect 50764 62972 50820 62974
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 49868 62412 49924 62468
rect 50092 62466 50148 62468
rect 50092 62414 50094 62466
rect 50094 62414 50146 62466
rect 50146 62414 50148 62466
rect 50092 62412 50148 62414
rect 48860 62188 48916 62244
rect 49308 62076 49364 62132
rect 51324 62524 51380 62580
rect 50428 62076 50484 62132
rect 51100 62076 51156 62132
rect 50428 61628 50484 61684
rect 50204 60786 50260 60788
rect 50204 60734 50206 60786
rect 50206 60734 50258 60786
rect 50258 60734 50260 60786
rect 50204 60732 50260 60734
rect 48524 59836 48580 59892
rect 48300 59612 48356 59668
rect 49196 60114 49252 60116
rect 49196 60062 49198 60114
rect 49198 60062 49250 60114
rect 49250 60062 49252 60114
rect 49196 60060 49252 60062
rect 48748 60002 48804 60004
rect 48748 59950 48750 60002
rect 48750 59950 48802 60002
rect 48802 59950 48804 60002
rect 48748 59948 48804 59950
rect 48972 59612 49028 59668
rect 48748 59218 48804 59220
rect 48748 59166 48750 59218
rect 48750 59166 48802 59218
rect 48802 59166 48804 59218
rect 48748 59164 48804 59166
rect 48412 56364 48468 56420
rect 48748 57538 48804 57540
rect 48748 57486 48750 57538
rect 48750 57486 48802 57538
rect 48802 57486 48804 57538
rect 48748 57484 48804 57486
rect 48524 56028 48580 56084
rect 48636 56140 48692 56196
rect 48300 55970 48356 55972
rect 48300 55918 48302 55970
rect 48302 55918 48354 55970
rect 48354 55918 48356 55970
rect 48300 55916 48356 55918
rect 47292 54684 47348 54740
rect 48300 55468 48356 55524
rect 47404 54514 47460 54516
rect 47404 54462 47406 54514
rect 47406 54462 47458 54514
rect 47458 54462 47460 54514
rect 47404 54460 47460 54462
rect 47404 53676 47460 53732
rect 47292 53506 47348 53508
rect 47292 53454 47294 53506
rect 47294 53454 47346 53506
rect 47346 53454 47348 53506
rect 47292 53452 47348 53454
rect 47180 53228 47236 53284
rect 47628 53340 47684 53396
rect 47068 52444 47124 52500
rect 46732 49644 46788 49700
rect 46508 49138 46564 49140
rect 46508 49086 46510 49138
rect 46510 49086 46562 49138
rect 46562 49086 46564 49138
rect 46508 49084 46564 49086
rect 46060 48914 46116 48916
rect 46060 48862 46062 48914
rect 46062 48862 46114 48914
rect 46114 48862 46116 48914
rect 46060 48860 46116 48862
rect 46956 51100 47012 51156
rect 46844 50204 46900 50260
rect 47068 50092 47124 50148
rect 47068 49810 47124 49812
rect 47068 49758 47070 49810
rect 47070 49758 47122 49810
rect 47122 49758 47124 49810
rect 47068 49756 47124 49758
rect 46284 48130 46340 48132
rect 46284 48078 46286 48130
rect 46286 48078 46338 48130
rect 46338 48078 46340 48130
rect 46284 48076 46340 48078
rect 47068 48748 47124 48804
rect 48188 55074 48244 55076
rect 48188 55022 48190 55074
rect 48190 55022 48242 55074
rect 48242 55022 48244 55074
rect 48188 55020 48244 55022
rect 47852 54908 47908 54964
rect 48188 54796 48244 54852
rect 47964 54348 48020 54404
rect 48188 53788 48244 53844
rect 48076 53228 48132 53284
rect 47740 52556 47796 52612
rect 47740 52108 47796 52164
rect 47964 52332 48020 52388
rect 48076 52668 48132 52724
rect 47852 52220 47908 52276
rect 47516 51490 47572 51492
rect 47516 51438 47518 51490
rect 47518 51438 47570 51490
rect 47570 51438 47572 51490
rect 47516 51436 47572 51438
rect 48076 52108 48132 52164
rect 48412 54124 48468 54180
rect 48412 53788 48468 53844
rect 48412 52444 48468 52500
rect 48412 52220 48468 52276
rect 48076 51212 48132 51268
rect 47404 50092 47460 50148
rect 47404 49922 47460 49924
rect 47404 49870 47406 49922
rect 47406 49870 47458 49922
rect 47458 49870 47460 49922
rect 47404 49868 47460 49870
rect 47404 48636 47460 48692
rect 47964 50316 48020 50372
rect 47852 49868 47908 49924
rect 47852 49138 47908 49140
rect 47852 49086 47854 49138
rect 47854 49086 47906 49138
rect 47906 49086 47908 49138
rect 47852 49084 47908 49086
rect 46844 47516 46900 47572
rect 46844 46898 46900 46900
rect 46844 46846 46846 46898
rect 46846 46846 46898 46898
rect 46898 46846 46900 46898
rect 46844 46844 46900 46846
rect 46956 45106 47012 45108
rect 46956 45054 46958 45106
rect 46958 45054 47010 45106
rect 47010 45054 47012 45106
rect 46956 45052 47012 45054
rect 47068 44044 47124 44100
rect 45948 36988 46004 37044
rect 46620 36988 46676 37044
rect 45052 34018 45108 34020
rect 45052 33966 45054 34018
rect 45054 33966 45106 34018
rect 45106 33966 45108 34018
rect 45052 33964 45108 33966
rect 46060 34188 46116 34244
rect 46396 33458 46452 33460
rect 46396 33406 46398 33458
rect 46398 33406 46450 33458
rect 46450 33406 46452 33458
rect 46396 33404 46452 33406
rect 45388 33180 45444 33236
rect 46620 33292 46676 33348
rect 46956 33234 47012 33236
rect 46956 33182 46958 33234
rect 46958 33182 47010 33234
rect 47010 33182 47012 33234
rect 46956 33180 47012 33182
rect 47964 48354 48020 48356
rect 47964 48302 47966 48354
rect 47966 48302 48018 48354
rect 48018 48302 48020 48354
rect 47964 48300 48020 48302
rect 48300 51266 48356 51268
rect 48300 51214 48302 51266
rect 48302 51214 48354 51266
rect 48354 51214 48356 51266
rect 48300 51212 48356 51214
rect 48300 50594 48356 50596
rect 48300 50542 48302 50594
rect 48302 50542 48354 50594
rect 48354 50542 48356 50594
rect 48300 50540 48356 50542
rect 48636 55468 48692 55524
rect 48860 56082 48916 56084
rect 48860 56030 48862 56082
rect 48862 56030 48914 56082
rect 48914 56030 48916 56082
rect 48860 56028 48916 56030
rect 49308 59276 49364 59332
rect 49420 59948 49476 60004
rect 49084 58546 49140 58548
rect 49084 58494 49086 58546
rect 49086 58494 49138 58546
rect 49138 58494 49140 58546
rect 49084 58492 49140 58494
rect 48972 55244 49028 55300
rect 48636 54460 48692 54516
rect 49196 55468 49252 55524
rect 49196 55298 49252 55300
rect 49196 55246 49198 55298
rect 49198 55246 49250 55298
rect 49250 55246 49252 55298
rect 49196 55244 49252 55246
rect 49084 54796 49140 54852
rect 49308 54908 49364 54964
rect 48860 54738 48916 54740
rect 48860 54686 48862 54738
rect 48862 54686 48914 54738
rect 48914 54686 48916 54738
rect 48860 54684 48916 54686
rect 48748 53842 48804 53844
rect 48748 53790 48750 53842
rect 48750 53790 48802 53842
rect 48802 53790 48804 53842
rect 48748 53788 48804 53790
rect 49196 53618 49252 53620
rect 49196 53566 49198 53618
rect 49198 53566 49250 53618
rect 49250 53566 49252 53618
rect 49196 53564 49252 53566
rect 48860 53452 48916 53508
rect 49084 53340 49140 53396
rect 48636 52444 48692 52500
rect 48636 52162 48692 52164
rect 48636 52110 48638 52162
rect 48638 52110 48690 52162
rect 48690 52110 48692 52162
rect 48636 52108 48692 52110
rect 49196 52386 49252 52388
rect 49196 52334 49198 52386
rect 49198 52334 49250 52386
rect 49250 52334 49252 52386
rect 49196 52332 49252 52334
rect 48748 51324 48804 51380
rect 49084 51436 49140 51492
rect 48748 50540 48804 50596
rect 48972 50988 49028 51044
rect 48076 47964 48132 48020
rect 48188 48076 48244 48132
rect 47628 47570 47684 47572
rect 47628 47518 47630 47570
rect 47630 47518 47682 47570
rect 47682 47518 47684 47570
rect 47628 47516 47684 47518
rect 47292 46844 47348 46900
rect 47628 46674 47684 46676
rect 47628 46622 47630 46674
rect 47630 46622 47682 46674
rect 47682 46622 47684 46674
rect 47628 46620 47684 46622
rect 47516 45106 47572 45108
rect 47516 45054 47518 45106
rect 47518 45054 47570 45106
rect 47570 45054 47572 45106
rect 47516 45052 47572 45054
rect 48524 49980 48580 50036
rect 48412 49698 48468 49700
rect 48412 49646 48414 49698
rect 48414 49646 48466 49698
rect 48466 49646 48468 49698
rect 48412 49644 48468 49646
rect 48748 50034 48804 50036
rect 48748 49982 48750 50034
rect 48750 49982 48802 50034
rect 48802 49982 48804 50034
rect 48748 49980 48804 49982
rect 48860 49868 48916 49924
rect 49084 50876 49140 50932
rect 48636 48076 48692 48132
rect 49308 50204 49364 50260
rect 49196 49644 49252 49700
rect 49308 49308 49364 49364
rect 50316 60674 50372 60676
rect 50316 60622 50318 60674
rect 50318 60622 50370 60674
rect 50370 60622 50372 60674
rect 50316 60620 50372 60622
rect 49644 59612 49700 59668
rect 49756 59164 49812 59220
rect 49644 58492 49700 58548
rect 49532 57762 49588 57764
rect 49532 57710 49534 57762
rect 49534 57710 49586 57762
rect 49586 57710 49588 57762
rect 49532 57708 49588 57710
rect 49644 56364 49700 56420
rect 49644 55522 49700 55524
rect 49644 55470 49646 55522
rect 49646 55470 49698 55522
rect 49698 55470 49700 55522
rect 49644 55468 49700 55470
rect 49868 57484 49924 57540
rect 50316 60002 50372 60004
rect 50316 59950 50318 60002
rect 50318 59950 50370 60002
rect 50370 59950 50372 60002
rect 50316 59948 50372 59950
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50204 59836 50260 59892
rect 51324 62188 51380 62244
rect 51212 61682 51268 61684
rect 51212 61630 51214 61682
rect 51214 61630 51266 61682
rect 51266 61630 51268 61682
rect 51212 61628 51268 61630
rect 51100 61068 51156 61124
rect 50876 59836 50932 59892
rect 50988 60732 51044 60788
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50988 59500 51044 59556
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50540 57538 50596 57540
rect 50540 57486 50542 57538
rect 50542 57486 50594 57538
rect 50594 57486 50596 57538
rect 50540 57484 50596 57486
rect 50428 56812 50484 56868
rect 49868 55692 49924 55748
rect 50204 56082 50260 56084
rect 50204 56030 50206 56082
rect 50206 56030 50258 56082
rect 50258 56030 50260 56082
rect 50204 56028 50260 56030
rect 50988 57538 51044 57540
rect 50988 57486 50990 57538
rect 50990 57486 51042 57538
rect 51042 57486 51044 57538
rect 50988 57484 51044 57486
rect 51324 59500 51380 59556
rect 51324 58044 51380 58100
rect 51548 60674 51604 60676
rect 51548 60622 51550 60674
rect 51550 60622 51602 60674
rect 51602 60622 51604 60674
rect 51548 60620 51604 60622
rect 52332 66162 52388 66164
rect 52332 66110 52334 66162
rect 52334 66110 52386 66162
rect 52386 66110 52388 66162
rect 52332 66108 52388 66110
rect 51996 65996 52052 66052
rect 53116 115948 53172 116004
rect 52668 67058 52724 67060
rect 52668 67006 52670 67058
rect 52670 67006 52722 67058
rect 52722 67006 52724 67058
rect 52668 67004 52724 67006
rect 52892 62354 52948 62356
rect 52892 62302 52894 62354
rect 52894 62302 52946 62354
rect 52946 62302 52948 62354
rect 52892 62300 52948 62302
rect 52444 61628 52500 61684
rect 52220 61346 52276 61348
rect 52220 61294 52222 61346
rect 52222 61294 52274 61346
rect 52274 61294 52276 61346
rect 52220 61292 52276 61294
rect 52668 61180 52724 61236
rect 52668 61010 52724 61012
rect 52668 60958 52670 61010
rect 52670 60958 52722 61010
rect 52722 60958 52724 61010
rect 52668 60956 52724 60958
rect 51884 60002 51940 60004
rect 51884 59950 51886 60002
rect 51886 59950 51938 60002
rect 51938 59950 51940 60002
rect 51884 59948 51940 59950
rect 51212 57484 51268 57540
rect 51772 59836 51828 59892
rect 50876 56588 50932 56644
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 51100 56194 51156 56196
rect 51100 56142 51102 56194
rect 51102 56142 51154 56194
rect 51154 56142 51156 56194
rect 51100 56140 51156 56142
rect 50652 56028 50708 56084
rect 50316 55580 50372 55636
rect 50540 55804 50596 55860
rect 50652 55580 50708 55636
rect 50092 55468 50148 55524
rect 50540 55298 50596 55300
rect 50540 55246 50542 55298
rect 50542 55246 50594 55298
rect 50594 55246 50596 55298
rect 50540 55244 50596 55246
rect 49756 54908 49812 54964
rect 50556 54906 50612 54908
rect 49532 54796 49588 54852
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50988 54908 51044 54964
rect 51212 54908 51268 54964
rect 49644 54572 49700 54628
rect 49868 54514 49924 54516
rect 49868 54462 49870 54514
rect 49870 54462 49922 54514
rect 49922 54462 49924 54514
rect 49868 54460 49924 54462
rect 50204 54514 50260 54516
rect 50204 54462 50206 54514
rect 50206 54462 50258 54514
rect 50258 54462 50260 54514
rect 50204 54460 50260 54462
rect 49644 53954 49700 53956
rect 49644 53902 49646 53954
rect 49646 53902 49698 53954
rect 49698 53902 49700 53954
rect 49644 53900 49700 53902
rect 49756 53788 49812 53844
rect 49644 52108 49700 52164
rect 49644 51602 49700 51604
rect 49644 51550 49646 51602
rect 49646 51550 49698 51602
rect 49698 51550 49700 51602
rect 49644 51548 49700 51550
rect 49420 50540 49476 50596
rect 49756 51212 49812 51268
rect 49532 49532 49588 49588
rect 49420 49084 49476 49140
rect 49308 49026 49364 49028
rect 49308 48974 49310 49026
rect 49310 48974 49362 49026
rect 49362 48974 49364 49026
rect 49308 48972 49364 48974
rect 49644 49026 49700 49028
rect 49644 48974 49646 49026
rect 49646 48974 49698 49026
rect 49698 48974 49700 49026
rect 49644 48972 49700 48974
rect 49756 49756 49812 49812
rect 48412 45612 48468 45668
rect 48972 46956 49028 47012
rect 48972 45612 49028 45668
rect 48636 45330 48692 45332
rect 48636 45278 48638 45330
rect 48638 45278 48690 45330
rect 48690 45278 48692 45330
rect 48636 45276 48692 45278
rect 47852 44044 47908 44100
rect 48076 44098 48132 44100
rect 48076 44046 48078 44098
rect 48078 44046 48130 44098
rect 48130 44046 48132 44098
rect 48076 44044 48132 44046
rect 48300 43426 48356 43428
rect 48300 43374 48302 43426
rect 48302 43374 48354 43426
rect 48354 43374 48356 43426
rect 48300 43372 48356 43374
rect 48188 42754 48244 42756
rect 48188 42702 48190 42754
rect 48190 42702 48242 42754
rect 48242 42702 48244 42754
rect 48188 42700 48244 42702
rect 47740 42530 47796 42532
rect 47740 42478 47742 42530
rect 47742 42478 47794 42530
rect 47794 42478 47796 42530
rect 47740 42476 47796 42478
rect 48300 41858 48356 41860
rect 48300 41806 48302 41858
rect 48302 41806 48354 41858
rect 48354 41806 48356 41858
rect 48300 41804 48356 41806
rect 47628 40908 47684 40964
rect 47404 40236 47460 40292
rect 47404 39452 47460 39508
rect 47180 34242 47236 34244
rect 47180 34190 47182 34242
rect 47182 34190 47234 34242
rect 47234 34190 47236 34242
rect 47180 34188 47236 34190
rect 44716 26962 44772 26964
rect 44716 26910 44718 26962
rect 44718 26910 44770 26962
rect 44770 26910 44772 26962
rect 44716 26908 44772 26910
rect 44716 23826 44772 23828
rect 44716 23774 44718 23826
rect 44718 23774 44770 23826
rect 44770 23774 44772 23826
rect 44716 23772 44772 23774
rect 44268 22092 44324 22148
rect 45052 21980 45108 22036
rect 44492 21698 44548 21700
rect 44492 21646 44494 21698
rect 44494 21646 44546 21698
rect 44546 21646 44548 21698
rect 44492 21644 44548 21646
rect 45052 21474 45108 21476
rect 45052 21422 45054 21474
rect 45054 21422 45106 21474
rect 45106 21422 45108 21474
rect 45052 21420 45108 21422
rect 43596 6636 43652 6692
rect 46060 27298 46116 27300
rect 46060 27246 46062 27298
rect 46062 27246 46114 27298
rect 46114 27246 46116 27298
rect 46060 27244 46116 27246
rect 46844 27132 46900 27188
rect 46620 26962 46676 26964
rect 46620 26910 46622 26962
rect 46622 26910 46674 26962
rect 46674 26910 46676 26962
rect 46620 26908 46676 26910
rect 46060 23938 46116 23940
rect 46060 23886 46062 23938
rect 46062 23886 46114 23938
rect 46114 23886 46116 23938
rect 46060 23884 46116 23886
rect 46620 23826 46676 23828
rect 46620 23774 46622 23826
rect 46622 23774 46674 23826
rect 46674 23774 46676 23826
rect 46620 23772 46676 23774
rect 46844 23660 46900 23716
rect 45500 21980 45556 22036
rect 47292 27244 47348 27300
rect 48412 39730 48468 39732
rect 48412 39678 48414 39730
rect 48414 39678 48466 39730
rect 48466 39678 48468 39730
rect 48412 39676 48468 39678
rect 47740 33458 47796 33460
rect 47740 33406 47742 33458
rect 47742 33406 47794 33458
rect 47794 33406 47796 33458
rect 47740 33404 47796 33406
rect 48188 33346 48244 33348
rect 48188 33294 48190 33346
rect 48190 33294 48242 33346
rect 48242 33294 48244 33346
rect 48188 33292 48244 33294
rect 48188 31948 48244 32004
rect 47740 28476 47796 28532
rect 49532 46956 49588 47012
rect 49196 45666 49252 45668
rect 49196 45614 49198 45666
rect 49198 45614 49250 45666
rect 49250 45614 49252 45666
rect 49196 45612 49252 45614
rect 49420 45330 49476 45332
rect 49420 45278 49422 45330
rect 49422 45278 49474 45330
rect 49474 45278 49476 45330
rect 49420 45276 49476 45278
rect 48860 43036 48916 43092
rect 49532 43596 49588 43652
rect 49532 43372 49588 43428
rect 48748 41692 48804 41748
rect 49196 40908 49252 40964
rect 49420 41132 49476 41188
rect 48748 40402 48804 40404
rect 48748 40350 48750 40402
rect 48750 40350 48802 40402
rect 48802 40350 48804 40402
rect 48748 40348 48804 40350
rect 49420 40348 49476 40404
rect 50652 53676 50708 53732
rect 50540 53618 50596 53620
rect 50540 53566 50542 53618
rect 50542 53566 50594 53618
rect 50594 53566 50596 53618
rect 50540 53564 50596 53566
rect 51212 54514 51268 54516
rect 51212 54462 51214 54514
rect 51214 54462 51266 54514
rect 51266 54462 51268 54514
rect 51212 54460 51268 54462
rect 50876 54402 50932 54404
rect 50876 54350 50878 54402
rect 50878 54350 50930 54402
rect 50930 54350 50932 54402
rect 50876 54348 50932 54350
rect 51436 57148 51492 57204
rect 51548 56588 51604 56644
rect 51548 55804 51604 55860
rect 51436 55692 51492 55748
rect 51548 54684 51604 54740
rect 50764 53564 50820 53620
rect 51436 54236 51492 54292
rect 50652 53452 50708 53508
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50428 52556 50484 52612
rect 49980 51884 50036 51940
rect 50316 51938 50372 51940
rect 50316 51886 50318 51938
rect 50318 51886 50370 51938
rect 50370 51886 50372 51938
rect 50316 51884 50372 51886
rect 50204 50482 50260 50484
rect 50204 50430 50206 50482
rect 50206 50430 50258 50482
rect 50258 50430 50260 50482
rect 50204 50428 50260 50430
rect 49980 49756 50036 49812
rect 50092 48972 50148 49028
rect 49868 48354 49924 48356
rect 49868 48302 49870 48354
rect 49870 48302 49922 48354
rect 49922 48302 49924 48354
rect 49868 48300 49924 48302
rect 49868 46844 49924 46900
rect 49868 46674 49924 46676
rect 49868 46622 49870 46674
rect 49870 46622 49922 46674
rect 49922 46622 49924 46674
rect 49868 46620 49924 46622
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50428 51548 50484 51604
rect 50988 53730 51044 53732
rect 50988 53678 50990 53730
rect 50990 53678 51042 53730
rect 51042 53678 51044 53730
rect 50988 53676 51044 53678
rect 51324 53452 51380 53508
rect 50988 51938 51044 51940
rect 50988 51886 50990 51938
rect 50990 51886 51042 51938
rect 51042 51886 51044 51938
rect 50988 51884 51044 51886
rect 51100 51660 51156 51716
rect 51548 54012 51604 54068
rect 51660 54908 51716 54964
rect 51436 51660 51492 51716
rect 51548 53788 51604 53844
rect 52892 60508 52948 60564
rect 52780 59890 52836 59892
rect 52780 59838 52782 59890
rect 52782 59838 52834 59890
rect 52834 59838 52836 59890
rect 52780 59836 52836 59838
rect 52332 59388 52388 59444
rect 53004 60396 53060 60452
rect 52220 58604 52276 58660
rect 52780 58940 52836 58996
rect 51996 58268 52052 58324
rect 52444 57874 52500 57876
rect 52444 57822 52446 57874
rect 52446 57822 52498 57874
rect 52498 57822 52500 57874
rect 52444 57820 52500 57822
rect 51996 57596 52052 57652
rect 52668 57484 52724 57540
rect 52444 57260 52500 57316
rect 52220 56642 52276 56644
rect 52220 56590 52222 56642
rect 52222 56590 52274 56642
rect 52274 56590 52276 56642
rect 52220 56588 52276 56590
rect 52332 56252 52388 56308
rect 52332 56082 52388 56084
rect 52332 56030 52334 56082
rect 52334 56030 52386 56082
rect 52386 56030 52388 56082
rect 52332 56028 52388 56030
rect 51996 55916 52052 55972
rect 51772 54796 51828 54852
rect 51884 55468 51940 55524
rect 51996 55356 52052 55412
rect 52332 55356 52388 55412
rect 52108 55020 52164 55076
rect 52220 54684 52276 54740
rect 52108 54124 52164 54180
rect 51884 54012 51940 54068
rect 51996 53676 52052 53732
rect 51660 53340 51716 53396
rect 51772 53618 51828 53620
rect 51772 53566 51774 53618
rect 51774 53566 51826 53618
rect 51826 53566 51828 53618
rect 51772 53564 51828 53566
rect 52892 57148 52948 57204
rect 52668 56866 52724 56868
rect 52668 56814 52670 56866
rect 52670 56814 52722 56866
rect 52722 56814 52724 56866
rect 52668 56812 52724 56814
rect 58156 116562 58212 116564
rect 58156 116510 58158 116562
rect 58158 116510 58210 116562
rect 58210 116510 58212 116562
rect 58156 116508 58212 116510
rect 56364 116060 56420 116116
rect 54460 113820 54516 113876
rect 56924 114770 56980 114772
rect 56924 114718 56926 114770
rect 56926 114718 56978 114770
rect 56978 114718 56980 114770
rect 56924 114716 56980 114718
rect 57484 114770 57540 114772
rect 57484 114718 57486 114770
rect 57486 114718 57538 114770
rect 57538 114718 57540 114770
rect 57484 114716 57540 114718
rect 59276 115836 59332 115892
rect 59500 116508 59556 116564
rect 56476 114658 56532 114660
rect 56476 114606 56478 114658
rect 56478 114606 56530 114658
rect 56530 114606 56532 114658
rect 56476 114604 56532 114606
rect 56924 102396 56980 102452
rect 55916 68796 55972 68852
rect 56476 68796 56532 68852
rect 54460 68236 54516 68292
rect 53228 68124 53284 68180
rect 53900 68012 53956 68068
rect 53340 65490 53396 65492
rect 53340 65438 53342 65490
rect 53342 65438 53394 65490
rect 53394 65438 53396 65490
rect 53340 65436 53396 65438
rect 54908 67116 54964 67172
rect 54796 66444 54852 66500
rect 54236 66220 54292 66276
rect 54012 66162 54068 66164
rect 54012 66110 54014 66162
rect 54014 66110 54066 66162
rect 54066 66110 54068 66162
rect 54012 66108 54068 66110
rect 53900 65436 53956 65492
rect 53676 64428 53732 64484
rect 54684 65884 54740 65940
rect 54908 65884 54964 65940
rect 54572 65436 54628 65492
rect 54236 65100 54292 65156
rect 54236 64482 54292 64484
rect 54236 64430 54238 64482
rect 54238 64430 54290 64482
rect 54290 64430 54292 64482
rect 54236 64428 54292 64430
rect 54012 64204 54068 64260
rect 53452 63308 53508 63364
rect 53340 62242 53396 62244
rect 53340 62190 53342 62242
rect 53342 62190 53394 62242
rect 53394 62190 53396 62242
rect 53340 62188 53396 62190
rect 53564 62524 53620 62580
rect 53788 61740 53844 61796
rect 53676 61180 53732 61236
rect 53564 60786 53620 60788
rect 53564 60734 53566 60786
rect 53566 60734 53618 60786
rect 53618 60734 53620 60786
rect 53564 60732 53620 60734
rect 54348 63868 54404 63924
rect 54348 63698 54404 63700
rect 54348 63646 54350 63698
rect 54350 63646 54402 63698
rect 54402 63646 54404 63698
rect 54348 63644 54404 63646
rect 55244 67004 55300 67060
rect 55692 67116 55748 67172
rect 55580 66946 55636 66948
rect 55580 66894 55582 66946
rect 55582 66894 55634 66946
rect 55634 66894 55636 66946
rect 55580 66892 55636 66894
rect 55356 66108 55412 66164
rect 55132 65660 55188 65716
rect 56252 67170 56308 67172
rect 56252 67118 56254 67170
rect 56254 67118 56306 67170
rect 56306 67118 56308 67170
rect 56252 67116 56308 67118
rect 56700 67564 56756 67620
rect 56140 66444 56196 66500
rect 56364 66892 56420 66948
rect 55916 66386 55972 66388
rect 55916 66334 55918 66386
rect 55918 66334 55970 66386
rect 55970 66334 55972 66386
rect 55916 66332 55972 66334
rect 55804 65996 55860 66052
rect 56588 66444 56644 66500
rect 56476 66050 56532 66052
rect 56476 65998 56478 66050
rect 56478 65998 56530 66050
rect 56530 65998 56532 66050
rect 56476 65996 56532 65998
rect 56364 65660 56420 65716
rect 56700 65884 56756 65940
rect 55916 65378 55972 65380
rect 55916 65326 55918 65378
rect 55918 65326 55970 65378
rect 55970 65326 55972 65378
rect 55916 65324 55972 65326
rect 55356 64706 55412 64708
rect 55356 64654 55358 64706
rect 55358 64654 55410 64706
rect 55410 64654 55412 64706
rect 55356 64652 55412 64654
rect 55916 64652 55972 64708
rect 55244 64204 55300 64260
rect 54796 62412 54852 62468
rect 55244 63644 55300 63700
rect 56700 65100 56756 65156
rect 56140 64652 56196 64708
rect 55356 63532 55412 63588
rect 56812 64092 56868 64148
rect 56140 63532 56196 63588
rect 56364 63532 56420 63588
rect 57932 92988 57988 93044
rect 57820 67618 57876 67620
rect 57820 67566 57822 67618
rect 57822 67566 57874 67618
rect 57874 67566 57876 67618
rect 57820 67564 57876 67566
rect 57596 67058 57652 67060
rect 57596 67006 57598 67058
rect 57598 67006 57650 67058
rect 57650 67006 57652 67058
rect 57596 67004 57652 67006
rect 57596 66274 57652 66276
rect 57596 66222 57598 66274
rect 57598 66222 57650 66274
rect 57650 66222 57652 66274
rect 57596 66220 57652 66222
rect 59948 116562 60004 116564
rect 59948 116510 59950 116562
rect 59950 116510 60002 116562
rect 60002 116510 60004 116562
rect 59948 116508 60004 116510
rect 60508 116508 60564 116564
rect 60060 115836 60116 115892
rect 58828 89516 58884 89572
rect 59276 68236 59332 68292
rect 58940 67116 58996 67172
rect 57932 66220 57988 66276
rect 55916 63084 55972 63140
rect 54460 62354 54516 62356
rect 54460 62302 54462 62354
rect 54462 62302 54514 62354
rect 54514 62302 54516 62354
rect 54460 62300 54516 62302
rect 55020 62354 55076 62356
rect 55020 62302 55022 62354
rect 55022 62302 55074 62354
rect 55074 62302 55076 62354
rect 55020 62300 55076 62302
rect 56252 62578 56308 62580
rect 56252 62526 56254 62578
rect 56254 62526 56306 62578
rect 56306 62526 56308 62578
rect 56252 62524 56308 62526
rect 55916 62300 55972 62356
rect 54124 61740 54180 61796
rect 55244 62188 55300 62244
rect 54124 61346 54180 61348
rect 54124 61294 54126 61346
rect 54126 61294 54178 61346
rect 54178 61294 54180 61346
rect 54124 61292 54180 61294
rect 53788 60956 53844 61012
rect 54348 61180 54404 61236
rect 55020 61180 55076 61236
rect 55020 60956 55076 61012
rect 54012 60562 54068 60564
rect 54012 60510 54014 60562
rect 54014 60510 54066 60562
rect 54066 60510 54068 60562
rect 54012 60508 54068 60510
rect 53900 60396 53956 60452
rect 53564 60002 53620 60004
rect 53564 59950 53566 60002
rect 53566 59950 53618 60002
rect 53618 59950 53620 60002
rect 53564 59948 53620 59950
rect 53340 56588 53396 56644
rect 53564 56812 53620 56868
rect 55020 60396 55076 60452
rect 55020 59948 55076 60004
rect 54908 59388 54964 59444
rect 55132 59836 55188 59892
rect 55468 62242 55524 62244
rect 55468 62190 55470 62242
rect 55470 62190 55522 62242
rect 55522 62190 55524 62242
rect 55468 62188 55524 62190
rect 55580 62076 55636 62132
rect 55356 60732 55412 60788
rect 56140 61964 56196 62020
rect 55804 61180 55860 61236
rect 56364 61180 56420 61236
rect 56364 60956 56420 61012
rect 56140 60732 56196 60788
rect 55356 60562 55412 60564
rect 55356 60510 55358 60562
rect 55358 60510 55410 60562
rect 55410 60510 55412 60562
rect 55356 60508 55412 60510
rect 55580 60002 55636 60004
rect 55580 59950 55582 60002
rect 55582 59950 55634 60002
rect 55634 59950 55636 60002
rect 55580 59948 55636 59950
rect 55468 59836 55524 59892
rect 54684 58994 54740 58996
rect 54684 58942 54686 58994
rect 54686 58942 54738 58994
rect 54738 58942 54740 58994
rect 54684 58940 54740 58942
rect 54460 58604 54516 58660
rect 54572 58716 54628 58772
rect 53788 58492 53844 58548
rect 54460 58322 54516 58324
rect 54460 58270 54462 58322
rect 54462 58270 54514 58322
rect 54514 58270 54516 58322
rect 54460 58268 54516 58270
rect 54236 57820 54292 57876
rect 53900 56866 53956 56868
rect 53900 56814 53902 56866
rect 53902 56814 53954 56866
rect 53954 56814 53956 56866
rect 53900 56812 53956 56814
rect 52556 55410 52612 55412
rect 52556 55358 52558 55410
rect 52558 55358 52610 55410
rect 52610 55358 52612 55410
rect 52556 55356 52612 55358
rect 52444 55020 52500 55076
rect 52332 53788 52388 53844
rect 51884 53058 51940 53060
rect 51884 53006 51886 53058
rect 51886 53006 51938 53058
rect 51938 53006 51940 53058
rect 51884 53004 51940 53006
rect 51772 52556 51828 52612
rect 51660 51548 51716 51604
rect 51996 52444 52052 52500
rect 50876 51436 50932 51492
rect 51436 51436 51492 51492
rect 50428 51212 50484 51268
rect 50540 51154 50596 51156
rect 50540 51102 50542 51154
rect 50542 51102 50594 51154
rect 50594 51102 50596 51154
rect 50540 51100 50596 51102
rect 50876 50988 50932 51044
rect 50876 50594 50932 50596
rect 50876 50542 50878 50594
rect 50878 50542 50930 50594
rect 50930 50542 50932 50594
rect 50876 50540 50932 50542
rect 51212 50594 51268 50596
rect 51212 50542 51214 50594
rect 51214 50542 51266 50594
rect 51266 50542 51268 50594
rect 51212 50540 51268 50542
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50988 50092 51044 50148
rect 50316 49138 50372 49140
rect 50316 49086 50318 49138
rect 50318 49086 50370 49138
rect 50370 49086 50372 49138
rect 50316 49084 50372 49086
rect 50204 48636 50260 48692
rect 50204 48076 50260 48132
rect 51324 49308 51380 49364
rect 50540 48860 50596 48916
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50764 48130 50820 48132
rect 50764 48078 50766 48130
rect 50766 48078 50818 48130
rect 50818 48078 50820 48130
rect 50764 48076 50820 48078
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50428 46844 50484 46900
rect 51548 50092 51604 50148
rect 51660 50316 51716 50372
rect 51548 49698 51604 49700
rect 51548 49646 51550 49698
rect 51550 49646 51602 49698
rect 51602 49646 51604 49698
rect 51548 49644 51604 49646
rect 51772 50204 51828 50260
rect 51884 49756 51940 49812
rect 51660 49196 51716 49252
rect 52220 52668 52276 52724
rect 52220 52386 52276 52388
rect 52220 52334 52222 52386
rect 52222 52334 52274 52386
rect 52274 52334 52276 52386
rect 52220 52332 52276 52334
rect 52892 55804 52948 55860
rect 53116 55468 53172 55524
rect 53452 55580 53508 55636
rect 53004 54738 53060 54740
rect 53004 54686 53006 54738
rect 53006 54686 53058 54738
rect 53058 54686 53060 54738
rect 53004 54684 53060 54686
rect 52780 53676 52836 53732
rect 53116 54012 53172 54068
rect 52892 53452 52948 53508
rect 52668 53228 52724 53284
rect 52780 52668 52836 52724
rect 53004 52444 53060 52500
rect 52444 51154 52500 51156
rect 52444 51102 52446 51154
rect 52446 51102 52498 51154
rect 52498 51102 52500 51154
rect 52444 51100 52500 51102
rect 52220 50988 52276 51044
rect 52108 49922 52164 49924
rect 52108 49870 52110 49922
rect 52110 49870 52162 49922
rect 52162 49870 52164 49922
rect 52108 49868 52164 49870
rect 52332 50204 52388 50260
rect 52108 49084 52164 49140
rect 52220 49196 52276 49252
rect 50316 46060 50372 46116
rect 49980 45612 50036 45668
rect 50204 45612 50260 45668
rect 49980 44322 50036 44324
rect 49980 44270 49982 44322
rect 49982 44270 50034 44322
rect 50034 44270 50036 44322
rect 49980 44268 50036 44270
rect 50652 46114 50708 46116
rect 50652 46062 50654 46114
rect 50654 46062 50706 46114
rect 50706 46062 50708 46114
rect 50652 46060 50708 46062
rect 50876 45724 50932 45780
rect 51436 45724 51492 45780
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50428 45276 50484 45332
rect 50540 44604 50596 44660
rect 51548 45500 51604 45556
rect 50988 45330 51044 45332
rect 50988 45278 50990 45330
rect 50990 45278 51042 45330
rect 51042 45278 51044 45330
rect 50988 45276 51044 45278
rect 51436 45330 51492 45332
rect 51436 45278 51438 45330
rect 51438 45278 51490 45330
rect 51490 45278 51492 45330
rect 51436 45276 51492 45278
rect 51772 45276 51828 45332
rect 50876 44604 50932 44660
rect 50428 44434 50484 44436
rect 50428 44382 50430 44434
rect 50430 44382 50482 44434
rect 50482 44382 50484 44434
rect 50428 44380 50484 44382
rect 50876 44098 50932 44100
rect 50876 44046 50878 44098
rect 50878 44046 50930 44098
rect 50930 44046 50932 44098
rect 50876 44044 50932 44046
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 49868 42754 49924 42756
rect 49868 42702 49870 42754
rect 49870 42702 49922 42754
rect 49922 42702 49924 42754
rect 49868 42700 49924 42702
rect 49756 42642 49812 42644
rect 49756 42590 49758 42642
rect 49758 42590 49810 42642
rect 49810 42590 49812 42642
rect 49756 42588 49812 42590
rect 49868 41804 49924 41860
rect 49868 41186 49924 41188
rect 49868 41134 49870 41186
rect 49870 41134 49922 41186
rect 49922 41134 49924 41186
rect 49868 41132 49924 41134
rect 49644 39676 49700 39732
rect 49868 39730 49924 39732
rect 49868 39678 49870 39730
rect 49870 39678 49922 39730
rect 49922 39678 49924 39730
rect 49868 39676 49924 39678
rect 48972 39506 49028 39508
rect 48972 39454 48974 39506
rect 48974 39454 49026 39506
rect 49026 39454 49028 39506
rect 48972 39452 49028 39454
rect 49196 39452 49252 39508
rect 48524 33404 48580 33460
rect 48412 31948 48468 32004
rect 48524 33180 48580 33236
rect 50204 39506 50260 39508
rect 50204 39454 50206 39506
rect 50206 39454 50258 39506
rect 50258 39454 50260 39506
rect 50204 39452 50260 39454
rect 48300 28476 48356 28532
rect 47852 27186 47908 27188
rect 47852 27134 47854 27186
rect 47854 27134 47906 27186
rect 47906 27134 47908 27186
rect 47852 27132 47908 27134
rect 47404 23826 47460 23828
rect 47404 23774 47406 23826
rect 47406 23774 47458 23826
rect 47458 23774 47460 23826
rect 47404 23772 47460 23774
rect 47180 22428 47236 22484
rect 46396 22204 46452 22260
rect 46844 22204 46900 22260
rect 46060 22146 46116 22148
rect 46060 22094 46062 22146
rect 46062 22094 46114 22146
rect 46114 22094 46116 22146
rect 46060 22092 46116 22094
rect 45836 20860 45892 20916
rect 45500 20130 45556 20132
rect 45500 20078 45502 20130
rect 45502 20078 45554 20130
rect 45554 20078 45556 20130
rect 45500 20076 45556 20078
rect 46620 20076 46676 20132
rect 46396 19794 46452 19796
rect 46396 19742 46398 19794
rect 46398 19742 46450 19794
rect 46450 19742 46452 19794
rect 46396 19740 46452 19742
rect 46060 6636 46116 6692
rect 43260 5234 43316 5236
rect 43260 5182 43262 5234
rect 43262 5182 43314 5234
rect 43314 5182 43316 5234
rect 43260 5180 43316 5182
rect 45948 4172 46004 4228
rect 46956 21980 47012 22036
rect 47180 21698 47236 21700
rect 47180 21646 47182 21698
rect 47182 21646 47234 21698
rect 47234 21646 47236 21698
rect 47180 21644 47236 21646
rect 46956 20130 47012 20132
rect 46956 20078 46958 20130
rect 46958 20078 47010 20130
rect 47010 20078 47012 20130
rect 46956 20076 47012 20078
rect 47180 20018 47236 20020
rect 47180 19966 47182 20018
rect 47182 19966 47234 20018
rect 47234 19966 47236 20018
rect 47180 19964 47236 19966
rect 48300 27132 48356 27188
rect 47852 23714 47908 23716
rect 47852 23662 47854 23714
rect 47854 23662 47906 23714
rect 47906 23662 47908 23714
rect 47852 23660 47908 23662
rect 47740 22258 47796 22260
rect 47740 22206 47742 22258
rect 47742 22206 47794 22258
rect 47794 22206 47796 22258
rect 47740 22204 47796 22206
rect 49420 28476 49476 28532
rect 48524 23660 48580 23716
rect 48188 22482 48244 22484
rect 48188 22430 48190 22482
rect 48190 22430 48242 22482
rect 48242 22430 48244 22482
rect 48188 22428 48244 22430
rect 48524 22428 48580 22484
rect 48524 22092 48580 22148
rect 47628 20914 47684 20916
rect 47628 20862 47630 20914
rect 47630 20862 47682 20914
rect 47682 20862 47684 20914
rect 47628 20860 47684 20862
rect 48300 20860 48356 20916
rect 48972 20914 49028 20916
rect 48972 20862 48974 20914
rect 48974 20862 49026 20914
rect 49026 20862 49028 20914
rect 48972 20860 49028 20862
rect 48300 20018 48356 20020
rect 48300 19966 48302 20018
rect 48302 19966 48354 20018
rect 48354 19966 48356 20018
rect 48300 19964 48356 19966
rect 47516 19740 47572 19796
rect 47740 19740 47796 19796
rect 44268 3442 44324 3444
rect 44268 3390 44270 3442
rect 44270 3390 44322 3442
rect 44322 3390 44324 3442
rect 44268 3388 44324 3390
rect 45164 3388 45220 3444
rect 48524 5180 48580 5236
rect 48076 4956 48132 5012
rect 48412 5010 48468 5012
rect 48412 4958 48414 5010
rect 48414 4958 48466 5010
rect 48466 4958 48468 5010
rect 48412 4956 48468 4958
rect 49196 5234 49252 5236
rect 49196 5182 49198 5234
rect 49198 5182 49250 5234
rect 49250 5182 49252 5234
rect 49196 5180 49252 5182
rect 49756 5180 49812 5236
rect 50764 43596 50820 43652
rect 50428 43036 50484 43092
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50876 41916 50932 41972
rect 51548 44492 51604 44548
rect 51324 44210 51380 44212
rect 51324 44158 51326 44210
rect 51326 44158 51378 44210
rect 51378 44158 51380 44210
rect 51324 44156 51380 44158
rect 51996 48802 52052 48804
rect 51996 48750 51998 48802
rect 51998 48750 52050 48802
rect 52050 48750 52052 48802
rect 51996 48748 52052 48750
rect 52220 46002 52276 46004
rect 52220 45950 52222 46002
rect 52222 45950 52274 46002
rect 52274 45950 52276 46002
rect 52220 45948 52276 45950
rect 52220 45612 52276 45668
rect 52444 48636 52500 48692
rect 51996 45218 52052 45220
rect 51996 45166 51998 45218
rect 51998 45166 52050 45218
rect 52050 45166 52052 45218
rect 51996 45164 52052 45166
rect 52668 50706 52724 50708
rect 52668 50654 52670 50706
rect 52670 50654 52722 50706
rect 52722 50654 52724 50706
rect 52668 50652 52724 50654
rect 53452 54012 53508 54068
rect 53228 52834 53284 52836
rect 53228 52782 53230 52834
rect 53230 52782 53282 52834
rect 53282 52782 53284 52834
rect 53228 52780 53284 52782
rect 53900 56364 53956 56420
rect 53788 56028 53844 56084
rect 53676 55970 53732 55972
rect 53676 55918 53678 55970
rect 53678 55918 53730 55970
rect 53730 55918 53732 55970
rect 53676 55916 53732 55918
rect 53788 55692 53844 55748
rect 53676 55298 53732 55300
rect 53676 55246 53678 55298
rect 53678 55246 53730 55298
rect 53730 55246 53732 55298
rect 53676 55244 53732 55246
rect 53900 55132 53956 55188
rect 54124 55410 54180 55412
rect 54124 55358 54126 55410
rect 54126 55358 54178 55410
rect 54178 55358 54180 55410
rect 54124 55356 54180 55358
rect 53564 53340 53620 53396
rect 53452 53228 53508 53284
rect 53340 51548 53396 51604
rect 52780 49698 52836 49700
rect 52780 49646 52782 49698
rect 52782 49646 52834 49698
rect 52834 49646 52836 49698
rect 52780 49644 52836 49646
rect 52668 49308 52724 49364
rect 52668 48860 52724 48916
rect 53004 48354 53060 48356
rect 53004 48302 53006 48354
rect 53006 48302 53058 48354
rect 53058 48302 53060 48354
rect 53004 48300 53060 48302
rect 52780 48188 52836 48244
rect 51548 42588 51604 42644
rect 51772 44156 51828 44212
rect 51772 42754 51828 42756
rect 51772 42702 51774 42754
rect 51774 42702 51826 42754
rect 51826 42702 51828 42754
rect 51772 42700 51828 42702
rect 51884 44044 51940 44100
rect 51436 42530 51492 42532
rect 51436 42478 51438 42530
rect 51438 42478 51490 42530
rect 51490 42478 51492 42530
rect 51436 42476 51492 42478
rect 50540 41074 50596 41076
rect 50540 41022 50542 41074
rect 50542 41022 50594 41074
rect 50594 41022 50596 41074
rect 50540 41020 50596 41022
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50988 41020 51044 41076
rect 51996 44380 52052 44436
rect 52444 44098 52500 44100
rect 52444 44046 52446 44098
rect 52446 44046 52498 44098
rect 52498 44046 52500 44098
rect 52444 44044 52500 44046
rect 53228 49308 53284 49364
rect 53676 52946 53732 52948
rect 53676 52894 53678 52946
rect 53678 52894 53730 52946
rect 53730 52894 53732 52946
rect 53676 52892 53732 52894
rect 53564 50988 53620 51044
rect 53676 52332 53732 52388
rect 54012 53116 54068 53172
rect 53900 51772 53956 51828
rect 54012 52556 54068 52612
rect 53900 51548 53956 51604
rect 54572 57820 54628 57876
rect 54348 57762 54404 57764
rect 54348 57710 54350 57762
rect 54350 57710 54402 57762
rect 54402 57710 54404 57762
rect 54348 57708 54404 57710
rect 54684 57372 54740 57428
rect 54460 56194 54516 56196
rect 54460 56142 54462 56194
rect 54462 56142 54514 56194
rect 54514 56142 54516 56194
rect 54460 56140 54516 56142
rect 55244 59164 55300 59220
rect 54684 55580 54740 55636
rect 54908 56082 54964 56084
rect 54908 56030 54910 56082
rect 54910 56030 54962 56082
rect 54962 56030 54964 56082
rect 54908 56028 54964 56030
rect 55356 58604 55412 58660
rect 55356 57484 55412 57540
rect 55468 57708 55524 57764
rect 55356 56364 55412 56420
rect 55132 55468 55188 55524
rect 54572 54514 54628 54516
rect 54572 54462 54574 54514
rect 54574 54462 54626 54514
rect 54626 54462 54628 54514
rect 54572 54460 54628 54462
rect 54348 54402 54404 54404
rect 54348 54350 54350 54402
rect 54350 54350 54402 54402
rect 54402 54350 54404 54402
rect 54348 54348 54404 54350
rect 54572 54236 54628 54292
rect 53788 50876 53844 50932
rect 53900 51212 53956 51268
rect 54348 53004 54404 53060
rect 53900 50652 53956 50708
rect 53788 50540 53844 50596
rect 53228 48076 53284 48132
rect 53452 46172 53508 46228
rect 53228 45164 53284 45220
rect 53228 44994 53284 44996
rect 53228 44942 53230 44994
rect 53230 44942 53282 44994
rect 53282 44942 53284 44994
rect 53228 44940 53284 44942
rect 53116 44156 53172 44212
rect 53676 49922 53732 49924
rect 53676 49870 53678 49922
rect 53678 49870 53730 49922
rect 53730 49870 53732 49922
rect 53676 49868 53732 49870
rect 54460 52162 54516 52164
rect 54460 52110 54462 52162
rect 54462 52110 54514 52162
rect 54514 52110 54516 52162
rect 54460 52108 54516 52110
rect 54012 49868 54068 49924
rect 53676 46508 53732 46564
rect 53676 45218 53732 45220
rect 53676 45166 53678 45218
rect 53678 45166 53730 45218
rect 53730 45166 53732 45218
rect 53676 45164 53732 45166
rect 54236 50652 54292 50708
rect 54684 53228 54740 53284
rect 54796 53004 54852 53060
rect 55244 52892 55300 52948
rect 54796 52332 54852 52388
rect 55580 57148 55636 57204
rect 55916 59218 55972 59220
rect 55916 59166 55918 59218
rect 55918 59166 55970 59218
rect 55970 59166 55972 59218
rect 55916 59164 55972 59166
rect 55804 58940 55860 58996
rect 56028 58322 56084 58324
rect 56028 58270 56030 58322
rect 56030 58270 56082 58322
rect 56082 58270 56084 58322
rect 56028 58268 56084 58270
rect 56252 59388 56308 59444
rect 56364 58716 56420 58772
rect 56700 62466 56756 62468
rect 56700 62414 56702 62466
rect 56702 62414 56754 62466
rect 56754 62414 56756 62466
rect 56700 62412 56756 62414
rect 56924 60620 56980 60676
rect 56812 59948 56868 60004
rect 56924 59836 56980 59892
rect 56924 59612 56980 59668
rect 57484 65378 57540 65380
rect 57484 65326 57486 65378
rect 57486 65326 57538 65378
rect 57538 65326 57540 65378
rect 57484 65324 57540 65326
rect 57372 65100 57428 65156
rect 57820 65324 57876 65380
rect 58044 65100 58100 65156
rect 57932 64764 57988 64820
rect 57484 64540 57540 64596
rect 59052 67004 59108 67060
rect 58716 66220 58772 66276
rect 58716 65548 58772 65604
rect 58828 64706 58884 64708
rect 58828 64654 58830 64706
rect 58830 64654 58882 64706
rect 58882 64654 58884 64706
rect 58828 64652 58884 64654
rect 58940 64594 58996 64596
rect 58940 64542 58942 64594
rect 58942 64542 58994 64594
rect 58994 64542 58996 64594
rect 58940 64540 58996 64542
rect 57820 64092 57876 64148
rect 57596 63922 57652 63924
rect 57596 63870 57598 63922
rect 57598 63870 57650 63922
rect 57650 63870 57652 63922
rect 57596 63868 57652 63870
rect 57372 63084 57428 63140
rect 57708 63308 57764 63364
rect 57260 60172 57316 60228
rect 57484 59948 57540 60004
rect 58268 63868 58324 63924
rect 58492 63868 58548 63924
rect 58044 62412 58100 62468
rect 58156 61404 58212 61460
rect 58044 60844 58100 60900
rect 57708 60674 57764 60676
rect 57708 60622 57710 60674
rect 57710 60622 57762 60674
rect 57762 60622 57764 60674
rect 57708 60620 57764 60622
rect 58156 60508 58212 60564
rect 57820 60002 57876 60004
rect 57820 59950 57822 60002
rect 57822 59950 57874 60002
rect 57874 59950 57876 60002
rect 57820 59948 57876 59950
rect 58940 63196 58996 63252
rect 58604 63138 58660 63140
rect 58604 63086 58606 63138
rect 58606 63086 58658 63138
rect 58658 63086 58660 63138
rect 58604 63084 58660 63086
rect 59164 63138 59220 63140
rect 59164 63086 59166 63138
rect 59166 63086 59218 63138
rect 59218 63086 59220 63138
rect 59164 63084 59220 63086
rect 58940 62466 58996 62468
rect 58940 62414 58942 62466
rect 58942 62414 58994 62466
rect 58994 62414 58996 62466
rect 58940 62412 58996 62414
rect 58380 60898 58436 60900
rect 58380 60846 58382 60898
rect 58382 60846 58434 60898
rect 58434 60846 58436 60898
rect 58380 60844 58436 60846
rect 58492 60786 58548 60788
rect 58492 60734 58494 60786
rect 58494 60734 58546 60786
rect 58546 60734 58548 60786
rect 58492 60732 58548 60734
rect 58604 60562 58660 60564
rect 58604 60510 58606 60562
rect 58606 60510 58658 60562
rect 58658 60510 58660 60562
rect 58604 60508 58660 60510
rect 59724 89570 59780 89572
rect 59724 89518 59726 89570
rect 59726 89518 59778 89570
rect 59778 89518 59780 89570
rect 59724 89516 59780 89518
rect 60732 89516 60788 89572
rect 59388 66386 59444 66388
rect 59388 66334 59390 66386
rect 59390 66334 59442 66386
rect 59442 66334 59444 66386
rect 59388 66332 59444 66334
rect 60620 67954 60676 67956
rect 60620 67902 60622 67954
rect 60622 67902 60674 67954
rect 60674 67902 60676 67954
rect 60620 67900 60676 67902
rect 60508 67564 60564 67620
rect 60508 66444 60564 66500
rect 60620 67004 60676 67060
rect 60172 64818 60228 64820
rect 60172 64766 60174 64818
rect 60174 64766 60226 64818
rect 60226 64766 60228 64818
rect 60172 64764 60228 64766
rect 60956 65378 61012 65380
rect 60956 65326 60958 65378
rect 60958 65326 61010 65378
rect 61010 65326 61012 65378
rect 60956 65324 61012 65326
rect 60620 64706 60676 64708
rect 60620 64654 60622 64706
rect 60622 64654 60674 64706
rect 60674 64654 60676 64706
rect 60620 64652 60676 64654
rect 59836 64540 59892 64596
rect 59724 64316 59780 64372
rect 58828 60844 58884 60900
rect 59500 64204 59556 64260
rect 59612 63138 59668 63140
rect 59612 63086 59614 63138
rect 59614 63086 59666 63138
rect 59666 63086 59668 63138
rect 59612 63084 59668 63086
rect 59836 64092 59892 64148
rect 59836 63922 59892 63924
rect 59836 63870 59838 63922
rect 59838 63870 59890 63922
rect 59890 63870 59892 63922
rect 59836 63868 59892 63870
rect 60956 63196 61012 63252
rect 60620 62412 60676 62468
rect 60284 61740 60340 61796
rect 59500 61628 59556 61684
rect 59612 60898 59668 60900
rect 59612 60846 59614 60898
rect 59614 60846 59666 60898
rect 59666 60846 59668 60898
rect 59612 60844 59668 60846
rect 59164 60786 59220 60788
rect 59164 60734 59166 60786
rect 59166 60734 59218 60786
rect 59218 60734 59220 60786
rect 59164 60732 59220 60734
rect 58940 60508 58996 60564
rect 59052 60620 59108 60676
rect 58716 60396 58772 60452
rect 58492 59948 58548 60004
rect 57148 59612 57204 59668
rect 57036 59388 57092 59444
rect 57820 59442 57876 59444
rect 57820 59390 57822 59442
rect 57822 59390 57874 59442
rect 57874 59390 57876 59442
rect 57820 59388 57876 59390
rect 56924 58940 56980 58996
rect 56700 58268 56756 58324
rect 56140 57820 56196 57876
rect 56028 57708 56084 57764
rect 55916 56924 55972 56980
rect 56140 56252 56196 56308
rect 56700 57874 56756 57876
rect 56700 57822 56702 57874
rect 56702 57822 56754 57874
rect 56754 57822 56756 57874
rect 56700 57820 56756 57822
rect 56700 56978 56756 56980
rect 56700 56926 56702 56978
rect 56702 56926 56754 56978
rect 56754 56926 56756 56978
rect 56700 56924 56756 56926
rect 55468 53452 55524 53508
rect 55692 54460 55748 54516
rect 56364 55970 56420 55972
rect 56364 55918 56366 55970
rect 56366 55918 56418 55970
rect 56418 55918 56420 55970
rect 56364 55916 56420 55918
rect 55804 55804 55860 55860
rect 54908 51772 54964 51828
rect 54908 51212 54964 51268
rect 54796 50764 54852 50820
rect 54572 50540 54628 50596
rect 54908 50652 54964 50708
rect 54236 49980 54292 50036
rect 54460 50092 54516 50148
rect 55020 50092 55076 50148
rect 54348 49922 54404 49924
rect 54348 49870 54350 49922
rect 54350 49870 54402 49922
rect 54402 49870 54404 49922
rect 54348 49868 54404 49870
rect 54236 49532 54292 49588
rect 56028 55804 56084 55860
rect 55916 54908 55972 54964
rect 55356 51436 55412 51492
rect 55468 51660 55524 51716
rect 55468 50988 55524 51044
rect 55356 50764 55412 50820
rect 55132 49868 55188 49924
rect 55244 49980 55300 50036
rect 54460 49084 54516 49140
rect 54684 49420 54740 49476
rect 54348 48972 54404 49028
rect 54012 48076 54068 48132
rect 54236 48076 54292 48132
rect 54572 47628 54628 47684
rect 55244 49026 55300 49028
rect 55244 48974 55246 49026
rect 55246 48974 55298 49026
rect 55298 48974 55300 49026
rect 55244 48972 55300 48974
rect 55692 51884 55748 51940
rect 55468 49980 55524 50036
rect 56364 55244 56420 55300
rect 56476 54460 56532 54516
rect 56252 53452 56308 53508
rect 54796 47964 54852 48020
rect 54684 46562 54740 46564
rect 54684 46510 54686 46562
rect 54686 46510 54738 46562
rect 54738 46510 54740 46562
rect 54684 46508 54740 46510
rect 53900 45948 53956 46004
rect 54124 45890 54180 45892
rect 54124 45838 54126 45890
rect 54126 45838 54178 45890
rect 54178 45838 54180 45890
rect 54124 45836 54180 45838
rect 53788 44940 53844 44996
rect 54012 45276 54068 45332
rect 53452 44098 53508 44100
rect 53452 44046 53454 44098
rect 53454 44046 53506 44098
rect 53506 44046 53508 44098
rect 53452 44044 53508 44046
rect 52892 43650 52948 43652
rect 52892 43598 52894 43650
rect 52894 43598 52946 43650
rect 52946 43598 52948 43650
rect 52892 43596 52948 43598
rect 53900 44210 53956 44212
rect 53900 44158 53902 44210
rect 53902 44158 53954 44210
rect 53954 44158 53956 44210
rect 53900 44156 53956 44158
rect 53788 43708 53844 43764
rect 54572 45276 54628 45332
rect 54460 44716 54516 44772
rect 54572 44828 54628 44884
rect 54124 44044 54180 44100
rect 54460 44156 54516 44212
rect 54236 43650 54292 43652
rect 54236 43598 54238 43650
rect 54238 43598 54290 43650
rect 54290 43598 54292 43650
rect 54236 43596 54292 43598
rect 53452 43148 53508 43204
rect 52220 42924 52276 42980
rect 53452 42812 53508 42868
rect 51884 41916 51940 41972
rect 51548 40460 51604 40516
rect 53676 42642 53732 42644
rect 53676 42590 53678 42642
rect 53678 42590 53730 42642
rect 53730 42590 53732 42642
rect 53676 42588 53732 42590
rect 52780 41858 52836 41860
rect 52780 41806 52782 41858
rect 52782 41806 52834 41858
rect 52834 41806 52836 41858
rect 52780 41804 52836 41806
rect 53452 41804 53508 41860
rect 52556 41692 52612 41748
rect 53900 41804 53956 41860
rect 53564 41244 53620 41300
rect 52668 41020 52724 41076
rect 53564 41020 53620 41076
rect 55244 48242 55300 48244
rect 55244 48190 55246 48242
rect 55246 48190 55298 48242
rect 55298 48190 55300 48242
rect 55244 48188 55300 48190
rect 55916 52386 55972 52388
rect 55916 52334 55918 52386
rect 55918 52334 55970 52386
rect 55970 52334 55972 52386
rect 55916 52332 55972 52334
rect 55020 46508 55076 46564
rect 55132 46396 55188 46452
rect 54236 41298 54292 41300
rect 54236 41246 54238 41298
rect 54238 41246 54290 41298
rect 54290 41246 54292 41298
rect 54236 41244 54292 41246
rect 53676 40514 53732 40516
rect 53676 40462 53678 40514
rect 53678 40462 53730 40514
rect 53730 40462 53732 40514
rect 53676 40460 53732 40462
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 53564 37436 53620 37492
rect 53564 36988 53620 37044
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 54236 37490 54292 37492
rect 54236 37438 54238 37490
rect 54238 37438 54290 37490
rect 54290 37438 54292 37490
rect 54236 37436 54292 37438
rect 54460 41804 54516 41860
rect 55356 46002 55412 46004
rect 55356 45950 55358 46002
rect 55358 45950 55410 46002
rect 55410 45950 55412 46002
rect 55356 45948 55412 45950
rect 55356 45612 55412 45668
rect 56252 51996 56308 52052
rect 56364 51884 56420 51940
rect 56476 51772 56532 51828
rect 56140 51436 56196 51492
rect 56476 50876 56532 50932
rect 56252 49644 56308 49700
rect 56364 49868 56420 49924
rect 56140 48130 56196 48132
rect 56140 48078 56142 48130
rect 56142 48078 56194 48130
rect 56194 48078 56196 48130
rect 56140 48076 56196 48078
rect 56140 47852 56196 47908
rect 55916 47458 55972 47460
rect 55916 47406 55918 47458
rect 55918 47406 55970 47458
rect 55970 47406 55972 47458
rect 55916 47404 55972 47406
rect 55692 45948 55748 46004
rect 55916 46396 55972 46452
rect 55356 44828 55412 44884
rect 55468 44940 55524 44996
rect 55244 44716 55300 44772
rect 54796 44044 54852 44100
rect 55356 43932 55412 43988
rect 55132 43596 55188 43652
rect 55244 43820 55300 43876
rect 54908 43372 54964 43428
rect 54908 42866 54964 42868
rect 54908 42814 54910 42866
rect 54910 42814 54962 42866
rect 54962 42814 54964 42866
rect 54908 42812 54964 42814
rect 55356 43708 55412 43764
rect 54572 37266 54628 37268
rect 54572 37214 54574 37266
rect 54574 37214 54626 37266
rect 54626 37214 54628 37266
rect 54572 37212 54628 37214
rect 53676 15202 53732 15204
rect 53676 15150 53678 15202
rect 53678 15150 53730 15202
rect 53730 15150 53732 15202
rect 53676 15148 53732 15150
rect 54684 37100 54740 37156
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 48524 3612 48580 3668
rect 49420 4562 49476 4564
rect 49420 4510 49422 4562
rect 49422 4510 49474 4562
rect 49474 4510 49476 4562
rect 49420 4508 49476 4510
rect 54460 15426 54516 15428
rect 54460 15374 54462 15426
rect 54462 15374 54514 15426
rect 54514 15374 54516 15426
rect 54460 15372 54516 15374
rect 54124 15148 54180 15204
rect 54012 4956 54068 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50316 4508 50372 4564
rect 51660 4508 51716 4564
rect 49532 3666 49588 3668
rect 49532 3614 49534 3666
rect 49534 3614 49586 3666
rect 49586 3614 49588 3666
rect 49532 3612 49588 3614
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 54460 4060 54516 4116
rect 54572 4172 54628 4228
rect 55132 37772 55188 37828
rect 55804 45164 55860 45220
rect 55916 44994 55972 44996
rect 55916 44942 55918 44994
rect 55918 44942 55970 44994
rect 55970 44942 55972 44994
rect 55916 44940 55972 44942
rect 55692 44716 55748 44772
rect 56476 49026 56532 49028
rect 56476 48974 56478 49026
rect 56478 48974 56530 49026
rect 56530 48974 56532 49026
rect 56476 48972 56532 48974
rect 56364 48748 56420 48804
rect 56364 47628 56420 47684
rect 56700 56252 56756 56308
rect 56700 54738 56756 54740
rect 56700 54686 56702 54738
rect 56702 54686 56754 54738
rect 56754 54686 56756 54738
rect 56700 54684 56756 54686
rect 57036 57708 57092 57764
rect 56924 54460 56980 54516
rect 57036 57484 57092 57540
rect 56924 53116 56980 53172
rect 56700 52668 56756 52724
rect 56812 52892 56868 52948
rect 56700 51436 56756 51492
rect 56924 51212 56980 51268
rect 57036 51996 57092 52052
rect 56812 50316 56868 50372
rect 56812 49532 56868 49588
rect 56924 48802 56980 48804
rect 56924 48750 56926 48802
rect 56926 48750 56978 48802
rect 56978 48750 56980 48802
rect 56924 48748 56980 48750
rect 56700 47628 56756 47684
rect 56812 48076 56868 48132
rect 56588 46396 56644 46452
rect 56364 45330 56420 45332
rect 56364 45278 56366 45330
rect 56366 45278 56418 45330
rect 56418 45278 56420 45330
rect 56364 45276 56420 45278
rect 55804 43932 55860 43988
rect 56364 43426 56420 43428
rect 56364 43374 56366 43426
rect 56366 43374 56418 43426
rect 56418 43374 56420 43426
rect 56364 43372 56420 43374
rect 56364 42866 56420 42868
rect 56364 42814 56366 42866
rect 56366 42814 56418 42866
rect 56418 42814 56420 42866
rect 56364 42812 56420 42814
rect 57036 48076 57092 48132
rect 57484 58716 57540 58772
rect 57596 58940 57652 58996
rect 57372 57708 57428 57764
rect 57260 56924 57316 56980
rect 57372 56252 57428 56308
rect 58492 59778 58548 59780
rect 58492 59726 58494 59778
rect 58494 59726 58546 59778
rect 58546 59726 58548 59778
rect 58492 59724 58548 59726
rect 58156 59612 58212 59668
rect 57820 57596 57876 57652
rect 57820 57148 57876 57204
rect 58492 59388 58548 59444
rect 59500 60786 59556 60788
rect 59500 60734 59502 60786
rect 59502 60734 59554 60786
rect 59554 60734 59556 60786
rect 59500 60732 59556 60734
rect 59948 60226 60004 60228
rect 59948 60174 59950 60226
rect 59950 60174 60002 60226
rect 60002 60174 60004 60226
rect 59948 60172 60004 60174
rect 59388 60002 59444 60004
rect 59388 59950 59390 60002
rect 59390 59950 59442 60002
rect 59442 59950 59444 60002
rect 59388 59948 59444 59950
rect 59724 60002 59780 60004
rect 59724 59950 59726 60002
rect 59726 59950 59778 60002
rect 59778 59950 59780 60002
rect 59724 59948 59780 59950
rect 60508 59948 60564 60004
rect 58604 58604 58660 58660
rect 58716 59052 58772 59108
rect 58268 58434 58324 58436
rect 58268 58382 58270 58434
rect 58270 58382 58322 58434
rect 58322 58382 58324 58434
rect 58268 58380 58324 58382
rect 58380 58156 58436 58212
rect 58380 57372 58436 57428
rect 58716 58268 58772 58324
rect 58156 56924 58212 56980
rect 57596 56082 57652 56084
rect 57596 56030 57598 56082
rect 57598 56030 57650 56082
rect 57650 56030 57652 56082
rect 57596 56028 57652 56030
rect 57484 55020 57540 55076
rect 57372 52834 57428 52836
rect 57372 52782 57374 52834
rect 57374 52782 57426 52834
rect 57426 52782 57428 52834
rect 57372 52780 57428 52782
rect 57596 54514 57652 54516
rect 57596 54462 57598 54514
rect 57598 54462 57650 54514
rect 57650 54462 57652 54514
rect 57596 54460 57652 54462
rect 59276 58716 59332 58772
rect 59164 58434 59220 58436
rect 59164 58382 59166 58434
rect 59166 58382 59218 58434
rect 59218 58382 59220 58434
rect 59164 58380 59220 58382
rect 58940 56978 58996 56980
rect 58940 56926 58942 56978
rect 58942 56926 58994 56978
rect 58994 56926 58996 56978
rect 58940 56924 58996 56926
rect 59388 58658 59444 58660
rect 59388 58606 59390 58658
rect 59390 58606 59442 58658
rect 59442 58606 59444 58658
rect 59388 58604 59444 58606
rect 60060 59724 60116 59780
rect 59612 58828 59668 58884
rect 60508 59500 60564 59556
rect 59948 58604 60004 58660
rect 59276 57596 59332 57652
rect 59500 57484 59556 57540
rect 59276 56978 59332 56980
rect 59276 56926 59278 56978
rect 59278 56926 59330 56978
rect 59330 56926 59332 56978
rect 59276 56924 59332 56926
rect 59836 56978 59892 56980
rect 59836 56926 59838 56978
rect 59838 56926 59890 56978
rect 59890 56926 59892 56978
rect 59836 56924 59892 56926
rect 59164 55858 59220 55860
rect 59164 55806 59166 55858
rect 59166 55806 59218 55858
rect 59218 55806 59220 55858
rect 59164 55804 59220 55806
rect 57932 55020 57988 55076
rect 58156 55074 58212 55076
rect 58156 55022 58158 55074
rect 58158 55022 58210 55074
rect 58210 55022 58212 55074
rect 58156 55020 58212 55022
rect 58940 55580 58996 55636
rect 58268 54908 58324 54964
rect 58604 55020 58660 55076
rect 57820 54684 57876 54740
rect 57820 54236 57876 54292
rect 58044 54460 58100 54516
rect 57932 53788 57988 53844
rect 57708 53116 57764 53172
rect 57820 53564 57876 53620
rect 57708 52834 57764 52836
rect 57708 52782 57710 52834
rect 57710 52782 57762 52834
rect 57762 52782 57764 52834
rect 57708 52780 57764 52782
rect 57260 52332 57316 52388
rect 57484 51490 57540 51492
rect 57484 51438 57486 51490
rect 57486 51438 57538 51490
rect 57538 51438 57540 51490
rect 57484 51436 57540 51438
rect 57708 51436 57764 51492
rect 57708 50764 57764 50820
rect 57484 49026 57540 49028
rect 57484 48974 57486 49026
rect 57486 48974 57538 49026
rect 57538 48974 57540 49026
rect 57484 48972 57540 48974
rect 57260 48188 57316 48244
rect 57484 48748 57540 48804
rect 57372 47458 57428 47460
rect 57372 47406 57374 47458
rect 57374 47406 57426 47458
rect 57426 47406 57428 47458
rect 57372 47404 57428 47406
rect 57596 48242 57652 48244
rect 57596 48190 57598 48242
rect 57598 48190 57650 48242
rect 57650 48190 57652 48242
rect 57596 48188 57652 48190
rect 58492 54514 58548 54516
rect 58492 54462 58494 54514
rect 58494 54462 58546 54514
rect 58546 54462 58548 54514
rect 58492 54460 58548 54462
rect 58492 53452 58548 53508
rect 58156 53228 58212 53284
rect 57708 47292 57764 47348
rect 57596 46956 57652 47012
rect 57260 45612 57316 45668
rect 57484 46508 57540 46564
rect 57596 45666 57652 45668
rect 57596 45614 57598 45666
rect 57598 45614 57650 45666
rect 57650 45614 57652 45666
rect 57596 45612 57652 45614
rect 57932 52556 57988 52612
rect 58044 52444 58100 52500
rect 58380 53116 58436 53172
rect 58828 54908 58884 54964
rect 59164 55298 59220 55300
rect 59164 55246 59166 55298
rect 59166 55246 59218 55298
rect 59218 55246 59220 55298
rect 59164 55244 59220 55246
rect 59500 56082 59556 56084
rect 59500 56030 59502 56082
rect 59502 56030 59554 56082
rect 59554 56030 59556 56082
rect 59500 56028 59556 56030
rect 59388 55410 59444 55412
rect 59388 55358 59390 55410
rect 59390 55358 59442 55410
rect 59442 55358 59444 55410
rect 59388 55356 59444 55358
rect 59500 55020 59556 55076
rect 60060 56642 60116 56644
rect 60060 56590 60062 56642
rect 60062 56590 60114 56642
rect 60114 56590 60116 56642
rect 60060 56588 60116 56590
rect 60620 57762 60676 57764
rect 60620 57710 60622 57762
rect 60622 57710 60674 57762
rect 60674 57710 60676 57762
rect 60620 57708 60676 57710
rect 60844 60508 60900 60564
rect 60956 60172 61012 60228
rect 60396 56812 60452 56868
rect 60508 57484 60564 57540
rect 60172 56028 60228 56084
rect 60172 55692 60228 55748
rect 58716 53564 58772 53620
rect 59052 54124 59108 54180
rect 58828 53116 58884 53172
rect 58716 52946 58772 52948
rect 58716 52894 58718 52946
rect 58718 52894 58770 52946
rect 58770 52894 58772 52946
rect 58716 52892 58772 52894
rect 58604 52556 58660 52612
rect 58380 52444 58436 52500
rect 59836 54124 59892 54180
rect 59612 53954 59668 53956
rect 59612 53902 59614 53954
rect 59614 53902 59666 53954
rect 59666 53902 59668 53954
rect 59612 53900 59668 53902
rect 59276 53842 59332 53844
rect 59276 53790 59278 53842
rect 59278 53790 59330 53842
rect 59330 53790 59332 53842
rect 59276 53788 59332 53790
rect 59836 53788 59892 53844
rect 59724 53676 59780 53732
rect 59388 53170 59444 53172
rect 59388 53118 59390 53170
rect 59390 53118 59442 53170
rect 59442 53118 59444 53170
rect 59388 53116 59444 53118
rect 59500 53004 59556 53060
rect 59276 52834 59332 52836
rect 59276 52782 59278 52834
rect 59278 52782 59330 52834
rect 59330 52782 59332 52834
rect 59276 52780 59332 52782
rect 58828 52332 58884 52388
rect 58828 51938 58884 51940
rect 58828 51886 58830 51938
rect 58830 51886 58882 51938
rect 58882 51886 58884 51938
rect 58828 51884 58884 51886
rect 58940 51772 58996 51828
rect 58604 51490 58660 51492
rect 58604 51438 58606 51490
rect 58606 51438 58658 51490
rect 58658 51438 58660 51490
rect 58604 51436 58660 51438
rect 58492 50764 58548 50820
rect 58828 50652 58884 50708
rect 58380 50316 58436 50372
rect 58828 50316 58884 50372
rect 58828 49420 58884 49476
rect 58716 48972 58772 49028
rect 59052 49644 59108 49700
rect 59164 51938 59220 51940
rect 59164 51886 59166 51938
rect 59166 51886 59218 51938
rect 59218 51886 59220 51938
rect 59164 51884 59220 51886
rect 59164 50876 59220 50932
rect 59388 52050 59444 52052
rect 59388 51998 59390 52050
rect 59390 51998 59442 52050
rect 59442 51998 59444 52050
rect 59388 51996 59444 51998
rect 59388 50706 59444 50708
rect 59388 50654 59390 50706
rect 59390 50654 59442 50706
rect 59442 50654 59444 50706
rect 59388 50652 59444 50654
rect 59724 51548 59780 51604
rect 60844 57484 60900 57540
rect 60732 56642 60788 56644
rect 60732 56590 60734 56642
rect 60734 56590 60786 56642
rect 60786 56590 60788 56642
rect 60732 56588 60788 56590
rect 61740 116508 61796 116564
rect 65916 116842 65972 116844
rect 65916 116790 65918 116842
rect 65918 116790 65970 116842
rect 65970 116790 65972 116842
rect 65916 116788 65972 116790
rect 66020 116842 66076 116844
rect 66020 116790 66022 116842
rect 66022 116790 66074 116842
rect 66074 116790 66076 116842
rect 66020 116788 66076 116790
rect 66124 116842 66180 116844
rect 66124 116790 66126 116842
rect 66126 116790 66178 116842
rect 66178 116790 66180 116842
rect 66124 116788 66180 116790
rect 65324 116508 65380 116564
rect 66444 116562 66500 116564
rect 66444 116510 66446 116562
rect 66446 116510 66498 116562
rect 66498 116510 66500 116562
rect 66444 116508 66500 116510
rect 62972 115724 63028 115780
rect 62972 114828 63028 114884
rect 61292 114604 61348 114660
rect 67340 116508 67396 116564
rect 69132 116562 69188 116564
rect 69132 116510 69134 116562
rect 69134 116510 69186 116562
rect 69186 116510 69188 116562
rect 69132 116508 69188 116510
rect 68796 115836 68852 115892
rect 69580 115890 69636 115892
rect 69580 115838 69582 115890
rect 69582 115838 69634 115890
rect 69634 115838 69636 115890
rect 69580 115836 69636 115838
rect 63644 114268 63700 114324
rect 64092 114322 64148 114324
rect 64092 114270 64094 114322
rect 64094 114270 64146 114322
rect 64146 114270 64148 114322
rect 64092 114268 64148 114270
rect 61292 94332 61348 94388
rect 61852 93548 61908 93604
rect 61964 86380 62020 86436
rect 62188 77756 62244 77812
rect 61404 67900 61460 67956
rect 61292 67058 61348 67060
rect 61292 67006 61294 67058
rect 61294 67006 61346 67058
rect 61346 67006 61348 67058
rect 61292 67004 61348 67006
rect 61180 63980 61236 64036
rect 61628 67900 61684 67956
rect 62188 68124 62244 68180
rect 62524 67730 62580 67732
rect 62524 67678 62526 67730
rect 62526 67678 62578 67730
rect 62578 67678 62580 67730
rect 62524 67676 62580 67678
rect 61516 65490 61572 65492
rect 61516 65438 61518 65490
rect 61518 65438 61570 65490
rect 61570 65438 61572 65490
rect 61516 65436 61572 65438
rect 61404 63026 61460 63028
rect 61404 62974 61406 63026
rect 61406 62974 61458 63026
rect 61458 62974 61460 63026
rect 61404 62972 61460 62974
rect 61180 61628 61236 61684
rect 61292 60786 61348 60788
rect 61292 60734 61294 60786
rect 61294 60734 61346 60786
rect 61346 60734 61348 60786
rect 61292 60732 61348 60734
rect 61292 60172 61348 60228
rect 61180 59218 61236 59220
rect 61180 59166 61182 59218
rect 61182 59166 61234 59218
rect 61234 59166 61236 59218
rect 61180 59164 61236 59166
rect 61516 62300 61572 62356
rect 61404 58380 61460 58436
rect 61404 58044 61460 58100
rect 61516 59612 61572 59668
rect 61404 56924 61460 56980
rect 62076 67004 62132 67060
rect 62636 66668 62692 66724
rect 62300 65602 62356 65604
rect 62300 65550 62302 65602
rect 62302 65550 62354 65602
rect 62354 65550 62356 65602
rect 62300 65548 62356 65550
rect 62412 65490 62468 65492
rect 62412 65438 62414 65490
rect 62414 65438 62466 65490
rect 62466 65438 62468 65490
rect 62412 65436 62468 65438
rect 61964 63980 62020 64036
rect 62972 67004 63028 67060
rect 63532 67116 63588 67172
rect 63980 67116 64036 67172
rect 63532 65884 63588 65940
rect 62076 63026 62132 63028
rect 62076 62974 62078 63026
rect 62078 62974 62130 63026
rect 62130 62974 62132 63026
rect 62076 62972 62132 62974
rect 61852 62354 61908 62356
rect 61852 62302 61854 62354
rect 61854 62302 61906 62354
rect 61906 62302 61908 62354
rect 61852 62300 61908 62302
rect 61852 60844 61908 60900
rect 61964 60786 62020 60788
rect 61964 60734 61966 60786
rect 61966 60734 62018 60786
rect 62018 60734 62020 60786
rect 61964 60732 62020 60734
rect 62636 64818 62692 64820
rect 62636 64766 62638 64818
rect 62638 64766 62690 64818
rect 62690 64766 62692 64818
rect 62636 64764 62692 64766
rect 62860 64428 62916 64484
rect 62636 63980 62692 64036
rect 62524 62524 62580 62580
rect 62412 60786 62468 60788
rect 62412 60734 62414 60786
rect 62414 60734 62466 60786
rect 62466 60734 62468 60786
rect 62412 60732 62468 60734
rect 61852 59388 61908 59444
rect 63196 65378 63252 65380
rect 63196 65326 63198 65378
rect 63198 65326 63250 65378
rect 63250 65326 63252 65378
rect 63196 65324 63252 65326
rect 64764 115500 64820 115556
rect 64428 114882 64484 114884
rect 64428 114830 64430 114882
rect 64430 114830 64482 114882
rect 64482 114830 64484 114882
rect 64428 114828 64484 114830
rect 65212 115500 65268 115556
rect 66332 115554 66388 115556
rect 66332 115502 66334 115554
rect 66334 115502 66386 115554
rect 66386 115502 66388 115554
rect 66332 115500 66388 115502
rect 67004 115500 67060 115556
rect 65916 115274 65972 115276
rect 65916 115222 65918 115274
rect 65918 115222 65970 115274
rect 65970 115222 65972 115274
rect 65916 115220 65972 115222
rect 66020 115274 66076 115276
rect 66020 115222 66022 115274
rect 66022 115222 66074 115274
rect 66074 115222 66076 115274
rect 66020 115220 66076 115222
rect 66124 115274 66180 115276
rect 66124 115222 66126 115274
rect 66126 115222 66178 115274
rect 66178 115222 66180 115274
rect 66124 115220 66180 115222
rect 70700 115612 70756 115668
rect 69020 115388 69076 115444
rect 69580 115388 69636 115444
rect 67004 114940 67060 114996
rect 65212 114268 65268 114324
rect 64092 67676 64148 67732
rect 64540 67116 64596 67172
rect 63980 65548 64036 65604
rect 64092 65996 64148 66052
rect 63868 65378 63924 65380
rect 63868 65326 63870 65378
rect 63870 65326 63922 65378
rect 63922 65326 63924 65378
rect 63868 65324 63924 65326
rect 63084 64204 63140 64260
rect 64540 65884 64596 65940
rect 64652 65996 64708 66052
rect 64988 65548 65044 65604
rect 63868 64428 63924 64484
rect 64092 64316 64148 64372
rect 63868 64092 63924 64148
rect 63756 63810 63812 63812
rect 63756 63758 63758 63810
rect 63758 63758 63810 63810
rect 63810 63758 63812 63810
rect 63756 63756 63812 63758
rect 62972 62914 63028 62916
rect 62972 62862 62974 62914
rect 62974 62862 63026 62914
rect 63026 62862 63028 62914
rect 62972 62860 63028 62862
rect 63084 62578 63140 62580
rect 63084 62526 63086 62578
rect 63086 62526 63138 62578
rect 63138 62526 63140 62578
rect 63084 62524 63140 62526
rect 63756 62860 63812 62916
rect 63980 63532 64036 63588
rect 64876 63980 64932 64036
rect 64204 63922 64260 63924
rect 64204 63870 64206 63922
rect 64206 63870 64258 63922
rect 64258 63870 64260 63922
rect 64204 63868 64260 63870
rect 64764 63756 64820 63812
rect 64764 62860 64820 62916
rect 63644 62354 63700 62356
rect 63644 62302 63646 62354
rect 63646 62302 63698 62354
rect 63698 62302 63700 62354
rect 63644 62300 63700 62302
rect 62636 59500 62692 59556
rect 61628 58716 61684 58772
rect 61628 57484 61684 57540
rect 60844 56082 60900 56084
rect 60844 56030 60846 56082
rect 60846 56030 60898 56082
rect 60898 56030 60900 56082
rect 60844 56028 60900 56030
rect 60620 54796 60676 54852
rect 60732 53900 60788 53956
rect 60508 53788 60564 53844
rect 60060 52556 60116 52612
rect 59948 51324 60004 51380
rect 59500 50428 59556 50484
rect 58940 48860 58996 48916
rect 58604 48748 58660 48804
rect 58156 48412 58212 48468
rect 58380 48130 58436 48132
rect 58380 48078 58382 48130
rect 58382 48078 58434 48130
rect 58434 48078 58436 48130
rect 58380 48076 58436 48078
rect 59500 50204 59556 50260
rect 58716 47628 58772 47684
rect 59612 47682 59668 47684
rect 59612 47630 59614 47682
rect 59614 47630 59666 47682
rect 59666 47630 59668 47682
rect 59612 47628 59668 47630
rect 59052 47458 59108 47460
rect 59052 47406 59054 47458
rect 59054 47406 59106 47458
rect 59106 47406 59108 47458
rect 59052 47404 59108 47406
rect 58268 47292 58324 47348
rect 58828 47346 58884 47348
rect 58828 47294 58830 47346
rect 58830 47294 58882 47346
rect 58882 47294 58884 47346
rect 58828 47292 58884 47294
rect 58716 46956 58772 47012
rect 57932 45836 57988 45892
rect 58156 46620 58212 46676
rect 57820 45276 57876 45332
rect 57148 45052 57204 45108
rect 55692 42588 55748 42644
rect 56812 42476 56868 42532
rect 56364 41916 56420 41972
rect 58604 46562 58660 46564
rect 58604 46510 58606 46562
rect 58606 46510 58658 46562
rect 58658 46510 58660 46562
rect 58604 46508 58660 46510
rect 59276 46508 59332 46564
rect 58604 45890 58660 45892
rect 58604 45838 58606 45890
rect 58606 45838 58658 45890
rect 58658 45838 58660 45890
rect 58604 45836 58660 45838
rect 58940 45890 58996 45892
rect 58940 45838 58942 45890
rect 58942 45838 58994 45890
rect 58994 45838 58996 45890
rect 58940 45836 58996 45838
rect 57820 43820 57876 43876
rect 57484 43650 57540 43652
rect 57484 43598 57486 43650
rect 57486 43598 57538 43650
rect 57538 43598 57540 43650
rect 57484 43596 57540 43598
rect 57932 42812 57988 42868
rect 58492 45106 58548 45108
rect 58492 45054 58494 45106
rect 58494 45054 58546 45106
rect 58546 45054 58548 45106
rect 58492 45052 58548 45054
rect 59276 45388 59332 45444
rect 58828 45218 58884 45220
rect 58828 45166 58830 45218
rect 58830 45166 58882 45218
rect 58882 45166 58884 45218
rect 58828 45164 58884 45166
rect 59388 45164 59444 45220
rect 58716 44940 58772 44996
rect 58380 44380 58436 44436
rect 58492 44828 58548 44884
rect 56364 40684 56420 40740
rect 55580 40236 55636 40292
rect 56476 40236 56532 40292
rect 56028 37772 56084 37828
rect 56364 37772 56420 37828
rect 56476 37212 56532 37268
rect 55468 37100 55524 37156
rect 54908 36988 54964 37044
rect 54796 5010 54852 5012
rect 54796 4958 54798 5010
rect 54798 4958 54850 5010
rect 54850 4958 54852 5010
rect 54796 4956 54852 4958
rect 58156 42530 58212 42532
rect 58156 42478 58158 42530
rect 58158 42478 58210 42530
rect 58210 42478 58212 42530
rect 58156 42476 58212 42478
rect 58156 42082 58212 42084
rect 58156 42030 58158 42082
rect 58158 42030 58210 42082
rect 58210 42030 58212 42082
rect 58156 42028 58212 42030
rect 57372 41132 57428 41188
rect 58268 41244 58324 41300
rect 58492 41132 58548 41188
rect 58940 45052 58996 45108
rect 57596 39564 57652 39620
rect 57708 40684 57764 40740
rect 57148 31052 57204 31108
rect 58156 40572 58212 40628
rect 59164 43260 59220 43316
rect 58716 42812 58772 42868
rect 59164 42028 59220 42084
rect 59612 45106 59668 45108
rect 59612 45054 59614 45106
rect 59614 45054 59666 45106
rect 59666 45054 59668 45106
rect 59612 45052 59668 45054
rect 59500 44828 59556 44884
rect 59500 44434 59556 44436
rect 59500 44382 59502 44434
rect 59502 44382 59554 44434
rect 59554 44382 59556 44434
rect 59500 44380 59556 44382
rect 59948 50594 60004 50596
rect 59948 50542 59950 50594
rect 59950 50542 60002 50594
rect 60002 50542 60004 50594
rect 59948 50540 60004 50542
rect 60060 48914 60116 48916
rect 60060 48862 60062 48914
rect 60062 48862 60114 48914
rect 60114 48862 60116 48914
rect 60060 48860 60116 48862
rect 59948 48748 60004 48804
rect 59836 47628 59892 47684
rect 61404 53676 61460 53732
rect 60508 53058 60564 53060
rect 60508 53006 60510 53058
rect 60510 53006 60562 53058
rect 60562 53006 60564 53058
rect 60508 53004 60564 53006
rect 62076 59218 62132 59220
rect 62076 59166 62078 59218
rect 62078 59166 62130 59218
rect 62130 59166 62132 59218
rect 62076 59164 62132 59166
rect 62188 58716 62244 58772
rect 62860 59442 62916 59444
rect 62860 59390 62862 59442
rect 62862 59390 62914 59442
rect 62914 59390 62916 59442
rect 62860 59388 62916 59390
rect 62748 59218 62804 59220
rect 62748 59166 62750 59218
rect 62750 59166 62802 59218
rect 62802 59166 62804 59218
rect 62748 59164 62804 59166
rect 62972 59052 63028 59108
rect 62860 58828 62916 58884
rect 62412 57820 62468 57876
rect 61964 57708 62020 57764
rect 61852 57538 61908 57540
rect 61852 57486 61854 57538
rect 61854 57486 61906 57538
rect 61906 57486 61908 57538
rect 61852 57484 61908 57486
rect 62300 56924 62356 56980
rect 62636 56978 62692 56980
rect 62636 56926 62638 56978
rect 62638 56926 62690 56978
rect 62690 56926 62692 56978
rect 62636 56924 62692 56926
rect 62524 56700 62580 56756
rect 62300 56476 62356 56532
rect 61740 55244 61796 55300
rect 61740 54236 61796 54292
rect 60284 52386 60340 52388
rect 60284 52334 60286 52386
rect 60286 52334 60338 52386
rect 60338 52334 60340 52386
rect 60284 52332 60340 52334
rect 60396 51772 60452 51828
rect 60284 51378 60340 51380
rect 60284 51326 60286 51378
rect 60286 51326 60338 51378
rect 60338 51326 60340 51378
rect 60284 51324 60340 51326
rect 60620 51324 60676 51380
rect 60620 49308 60676 49364
rect 60284 49084 60340 49140
rect 60732 48972 60788 49028
rect 60620 48748 60676 48804
rect 60396 48130 60452 48132
rect 60396 48078 60398 48130
rect 60398 48078 60450 48130
rect 60450 48078 60452 48130
rect 60396 48076 60452 48078
rect 60396 47628 60452 47684
rect 60284 45388 60340 45444
rect 60060 44828 60116 44884
rect 60060 44044 60116 44100
rect 59388 43596 59444 43652
rect 59612 43484 59668 43540
rect 59388 42588 59444 42644
rect 59388 42028 59444 42084
rect 59612 42476 59668 42532
rect 60284 43708 60340 43764
rect 59948 43314 60004 43316
rect 59948 43262 59950 43314
rect 59950 43262 60002 43314
rect 60002 43262 60004 43314
rect 59948 43260 60004 43262
rect 60060 43036 60116 43092
rect 59948 42812 60004 42868
rect 59836 41916 59892 41972
rect 59500 41298 59556 41300
rect 59500 41246 59502 41298
rect 59502 41246 59554 41298
rect 59554 41246 59556 41298
rect 59500 41244 59556 41246
rect 59052 41186 59108 41188
rect 59052 41134 59054 41186
rect 59054 41134 59106 41186
rect 59106 41134 59108 41186
rect 59052 41132 59108 41134
rect 58828 40572 58884 40628
rect 58604 40236 58660 40292
rect 58604 34690 58660 34692
rect 58604 34638 58606 34690
rect 58606 34638 58658 34690
rect 58658 34638 58660 34690
rect 58604 34636 58660 34638
rect 56364 9212 56420 9268
rect 58828 31948 58884 32004
rect 59836 22204 59892 22260
rect 55244 5010 55300 5012
rect 55244 4958 55246 5010
rect 55246 4958 55298 5010
rect 55298 4958 55300 5010
rect 55244 4956 55300 4958
rect 61404 52946 61460 52948
rect 61404 52894 61406 52946
rect 61406 52894 61458 52946
rect 61458 52894 61460 52946
rect 61404 52892 61460 52894
rect 60956 52332 61012 52388
rect 61516 52332 61572 52388
rect 61292 49644 61348 49700
rect 60844 46732 60900 46788
rect 61068 49420 61124 49476
rect 60844 46172 60900 46228
rect 60508 43484 60564 43540
rect 61180 48860 61236 48916
rect 61628 50652 61684 50708
rect 61628 50482 61684 50484
rect 61628 50430 61630 50482
rect 61630 50430 61682 50482
rect 61682 50430 61684 50482
rect 61628 50428 61684 50430
rect 61516 49308 61572 49364
rect 61852 53228 61908 53284
rect 61852 52444 61908 52500
rect 61740 49084 61796 49140
rect 61628 49026 61684 49028
rect 61628 48974 61630 49026
rect 61630 48974 61682 49026
rect 61682 48974 61684 49026
rect 61628 48972 61684 48974
rect 61516 48242 61572 48244
rect 61516 48190 61518 48242
rect 61518 48190 61570 48242
rect 61570 48190 61572 48242
rect 61516 48188 61572 48190
rect 61404 48130 61460 48132
rect 61404 48078 61406 48130
rect 61406 48078 61458 48130
rect 61458 48078 61460 48130
rect 61404 48076 61460 48078
rect 61292 47852 61348 47908
rect 61740 48354 61796 48356
rect 61740 48302 61742 48354
rect 61742 48302 61794 48354
rect 61794 48302 61796 48354
rect 61740 48300 61796 48302
rect 61852 48076 61908 48132
rect 61852 47852 61908 47908
rect 61404 45276 61460 45332
rect 61068 44604 61124 44660
rect 61292 45052 61348 45108
rect 62412 56306 62468 56308
rect 62412 56254 62414 56306
rect 62414 56254 62466 56306
rect 62466 56254 62468 56306
rect 62412 56252 62468 56254
rect 62076 55410 62132 55412
rect 62076 55358 62078 55410
rect 62078 55358 62130 55410
rect 62130 55358 62132 55410
rect 62076 55356 62132 55358
rect 62300 55298 62356 55300
rect 62300 55246 62302 55298
rect 62302 55246 62354 55298
rect 62354 55246 62356 55298
rect 62300 55244 62356 55246
rect 62300 55074 62356 55076
rect 62300 55022 62302 55074
rect 62302 55022 62354 55074
rect 62354 55022 62356 55074
rect 62300 55020 62356 55022
rect 62188 53618 62244 53620
rect 62188 53566 62190 53618
rect 62190 53566 62242 53618
rect 62242 53566 62244 53618
rect 62188 53564 62244 53566
rect 62076 53116 62132 53172
rect 62076 52780 62132 52836
rect 63308 56924 63364 56980
rect 62860 55970 62916 55972
rect 62860 55918 62862 55970
rect 62862 55918 62914 55970
rect 62914 55918 62916 55970
rect 62860 55916 62916 55918
rect 62860 55298 62916 55300
rect 62860 55246 62862 55298
rect 62862 55246 62914 55298
rect 62914 55246 62916 55298
rect 62860 55244 62916 55246
rect 62972 55186 63028 55188
rect 62972 55134 62974 55186
rect 62974 55134 63026 55186
rect 63026 55134 63028 55186
rect 62972 55132 63028 55134
rect 62860 54908 62916 54964
rect 63196 54572 63252 54628
rect 62748 54348 62804 54404
rect 62972 54402 63028 54404
rect 62972 54350 62974 54402
rect 62974 54350 63026 54402
rect 63026 54350 63028 54402
rect 62972 54348 63028 54350
rect 62524 53452 62580 53508
rect 62524 52444 62580 52500
rect 62636 53730 62692 53732
rect 62636 53678 62638 53730
rect 62638 53678 62690 53730
rect 62690 53678 62692 53730
rect 62636 53676 62692 53678
rect 62300 51996 62356 52052
rect 62412 52386 62468 52388
rect 62412 52334 62414 52386
rect 62414 52334 62466 52386
rect 62466 52334 62468 52386
rect 62412 52332 62468 52334
rect 62188 51884 62244 51940
rect 62076 50764 62132 50820
rect 62188 50594 62244 50596
rect 62188 50542 62190 50594
rect 62190 50542 62242 50594
rect 62242 50542 62244 50594
rect 62188 50540 62244 50542
rect 63084 52556 63140 52612
rect 62636 51324 62692 51380
rect 63084 51884 63140 51940
rect 62860 49644 62916 49700
rect 62412 48860 62468 48916
rect 62524 48188 62580 48244
rect 62524 47740 62580 47796
rect 62972 49138 63028 49140
rect 62972 49086 62974 49138
rect 62974 49086 63026 49138
rect 63026 49086 63028 49138
rect 62972 49084 63028 49086
rect 63308 53730 63364 53732
rect 63308 53678 63310 53730
rect 63310 53678 63362 53730
rect 63362 53678 63364 53730
rect 63308 53676 63364 53678
rect 63308 52834 63364 52836
rect 63308 52782 63310 52834
rect 63310 52782 63362 52834
rect 63362 52782 63364 52834
rect 63308 52780 63364 52782
rect 63532 60114 63588 60116
rect 63532 60062 63534 60114
rect 63534 60062 63586 60114
rect 63586 60062 63588 60114
rect 63532 60060 63588 60062
rect 63644 60508 63700 60564
rect 65916 113706 65972 113708
rect 65916 113654 65918 113706
rect 65918 113654 65970 113706
rect 65970 113654 65972 113706
rect 65916 113652 65972 113654
rect 66020 113706 66076 113708
rect 66020 113654 66022 113706
rect 66022 113654 66074 113706
rect 66074 113654 66076 113706
rect 66020 113652 66076 113654
rect 66124 113706 66180 113708
rect 66124 113654 66126 113706
rect 66126 113654 66178 113706
rect 66178 113654 66180 113706
rect 66124 113652 66180 113654
rect 67788 113372 67844 113428
rect 65916 112138 65972 112140
rect 65916 112086 65918 112138
rect 65918 112086 65970 112138
rect 65970 112086 65972 112138
rect 65916 112084 65972 112086
rect 66020 112138 66076 112140
rect 66020 112086 66022 112138
rect 66022 112086 66074 112138
rect 66074 112086 66076 112138
rect 66020 112084 66076 112086
rect 66124 112138 66180 112140
rect 66124 112086 66126 112138
rect 66126 112086 66178 112138
rect 66178 112086 66180 112138
rect 66124 112084 66180 112086
rect 65916 110570 65972 110572
rect 65916 110518 65918 110570
rect 65918 110518 65970 110570
rect 65970 110518 65972 110570
rect 65916 110516 65972 110518
rect 66020 110570 66076 110572
rect 66020 110518 66022 110570
rect 66022 110518 66074 110570
rect 66074 110518 66076 110570
rect 66020 110516 66076 110518
rect 66124 110570 66180 110572
rect 66124 110518 66126 110570
rect 66126 110518 66178 110570
rect 66178 110518 66180 110570
rect 66124 110516 66180 110518
rect 65916 109002 65972 109004
rect 65916 108950 65918 109002
rect 65918 108950 65970 109002
rect 65970 108950 65972 109002
rect 65916 108948 65972 108950
rect 66020 109002 66076 109004
rect 66020 108950 66022 109002
rect 66022 108950 66074 109002
rect 66074 108950 66076 109002
rect 66020 108948 66076 108950
rect 66124 109002 66180 109004
rect 66124 108950 66126 109002
rect 66126 108950 66178 109002
rect 66178 108950 66180 109002
rect 66124 108948 66180 108950
rect 65916 107434 65972 107436
rect 65916 107382 65918 107434
rect 65918 107382 65970 107434
rect 65970 107382 65972 107434
rect 65916 107380 65972 107382
rect 66020 107434 66076 107436
rect 66020 107382 66022 107434
rect 66022 107382 66074 107434
rect 66074 107382 66076 107434
rect 66020 107380 66076 107382
rect 66124 107434 66180 107436
rect 66124 107382 66126 107434
rect 66126 107382 66178 107434
rect 66178 107382 66180 107434
rect 66124 107380 66180 107382
rect 65916 105866 65972 105868
rect 65916 105814 65918 105866
rect 65918 105814 65970 105866
rect 65970 105814 65972 105866
rect 65916 105812 65972 105814
rect 66020 105866 66076 105868
rect 66020 105814 66022 105866
rect 66022 105814 66074 105866
rect 66074 105814 66076 105866
rect 66020 105812 66076 105814
rect 66124 105866 66180 105868
rect 66124 105814 66126 105866
rect 66126 105814 66178 105866
rect 66178 105814 66180 105866
rect 66124 105812 66180 105814
rect 65916 104298 65972 104300
rect 65916 104246 65918 104298
rect 65918 104246 65970 104298
rect 65970 104246 65972 104298
rect 65916 104244 65972 104246
rect 66020 104298 66076 104300
rect 66020 104246 66022 104298
rect 66022 104246 66074 104298
rect 66074 104246 66076 104298
rect 66020 104244 66076 104246
rect 66124 104298 66180 104300
rect 66124 104246 66126 104298
rect 66126 104246 66178 104298
rect 66178 104246 66180 104298
rect 66124 104244 66180 104246
rect 65916 102730 65972 102732
rect 65916 102678 65918 102730
rect 65918 102678 65970 102730
rect 65970 102678 65972 102730
rect 65916 102676 65972 102678
rect 66020 102730 66076 102732
rect 66020 102678 66022 102730
rect 66022 102678 66074 102730
rect 66074 102678 66076 102730
rect 66020 102676 66076 102678
rect 66124 102730 66180 102732
rect 66124 102678 66126 102730
rect 66126 102678 66178 102730
rect 66178 102678 66180 102730
rect 66124 102676 66180 102678
rect 65916 101162 65972 101164
rect 65916 101110 65918 101162
rect 65918 101110 65970 101162
rect 65970 101110 65972 101162
rect 65916 101108 65972 101110
rect 66020 101162 66076 101164
rect 66020 101110 66022 101162
rect 66022 101110 66074 101162
rect 66074 101110 66076 101162
rect 66020 101108 66076 101110
rect 66124 101162 66180 101164
rect 66124 101110 66126 101162
rect 66126 101110 66178 101162
rect 66178 101110 66180 101162
rect 66124 101108 66180 101110
rect 65916 99594 65972 99596
rect 65916 99542 65918 99594
rect 65918 99542 65970 99594
rect 65970 99542 65972 99594
rect 65916 99540 65972 99542
rect 66020 99594 66076 99596
rect 66020 99542 66022 99594
rect 66022 99542 66074 99594
rect 66074 99542 66076 99594
rect 66020 99540 66076 99542
rect 66124 99594 66180 99596
rect 66124 99542 66126 99594
rect 66126 99542 66178 99594
rect 66178 99542 66180 99594
rect 66124 99540 66180 99542
rect 65916 98026 65972 98028
rect 65916 97974 65918 98026
rect 65918 97974 65970 98026
rect 65970 97974 65972 98026
rect 65916 97972 65972 97974
rect 66020 98026 66076 98028
rect 66020 97974 66022 98026
rect 66022 97974 66074 98026
rect 66074 97974 66076 98026
rect 66020 97972 66076 97974
rect 66124 98026 66180 98028
rect 66124 97974 66126 98026
rect 66126 97974 66178 98026
rect 66178 97974 66180 98026
rect 66124 97972 66180 97974
rect 65916 96458 65972 96460
rect 65916 96406 65918 96458
rect 65918 96406 65970 96458
rect 65970 96406 65972 96458
rect 65916 96404 65972 96406
rect 66020 96458 66076 96460
rect 66020 96406 66022 96458
rect 66022 96406 66074 96458
rect 66074 96406 66076 96458
rect 66020 96404 66076 96406
rect 66124 96458 66180 96460
rect 66124 96406 66126 96458
rect 66126 96406 66178 96458
rect 66178 96406 66180 96458
rect 66124 96404 66180 96406
rect 65916 94890 65972 94892
rect 65916 94838 65918 94890
rect 65918 94838 65970 94890
rect 65970 94838 65972 94890
rect 65916 94836 65972 94838
rect 66020 94890 66076 94892
rect 66020 94838 66022 94890
rect 66022 94838 66074 94890
rect 66074 94838 66076 94890
rect 66020 94836 66076 94838
rect 66124 94890 66180 94892
rect 66124 94838 66126 94890
rect 66126 94838 66178 94890
rect 66178 94838 66180 94890
rect 66124 94836 66180 94838
rect 65916 93322 65972 93324
rect 65916 93270 65918 93322
rect 65918 93270 65970 93322
rect 65970 93270 65972 93322
rect 65916 93268 65972 93270
rect 66020 93322 66076 93324
rect 66020 93270 66022 93322
rect 66022 93270 66074 93322
rect 66074 93270 66076 93322
rect 66020 93268 66076 93270
rect 66124 93322 66180 93324
rect 66124 93270 66126 93322
rect 66126 93270 66178 93322
rect 66178 93270 66180 93322
rect 66124 93268 66180 93270
rect 65916 91754 65972 91756
rect 65916 91702 65918 91754
rect 65918 91702 65970 91754
rect 65970 91702 65972 91754
rect 65916 91700 65972 91702
rect 66020 91754 66076 91756
rect 66020 91702 66022 91754
rect 66022 91702 66074 91754
rect 66074 91702 66076 91754
rect 66020 91700 66076 91702
rect 66124 91754 66180 91756
rect 66124 91702 66126 91754
rect 66126 91702 66178 91754
rect 66178 91702 66180 91754
rect 66124 91700 66180 91702
rect 65916 90186 65972 90188
rect 65916 90134 65918 90186
rect 65918 90134 65970 90186
rect 65970 90134 65972 90186
rect 65916 90132 65972 90134
rect 66020 90186 66076 90188
rect 66020 90134 66022 90186
rect 66022 90134 66074 90186
rect 66074 90134 66076 90186
rect 66020 90132 66076 90134
rect 66124 90186 66180 90188
rect 66124 90134 66126 90186
rect 66126 90134 66178 90186
rect 66178 90134 66180 90186
rect 66124 90132 66180 90134
rect 65916 88618 65972 88620
rect 65916 88566 65918 88618
rect 65918 88566 65970 88618
rect 65970 88566 65972 88618
rect 65916 88564 65972 88566
rect 66020 88618 66076 88620
rect 66020 88566 66022 88618
rect 66022 88566 66074 88618
rect 66074 88566 66076 88618
rect 66020 88564 66076 88566
rect 66124 88618 66180 88620
rect 66124 88566 66126 88618
rect 66126 88566 66178 88618
rect 66178 88566 66180 88618
rect 66124 88564 66180 88566
rect 65916 87050 65972 87052
rect 65916 86998 65918 87050
rect 65918 86998 65970 87050
rect 65970 86998 65972 87050
rect 65916 86996 65972 86998
rect 66020 87050 66076 87052
rect 66020 86998 66022 87050
rect 66022 86998 66074 87050
rect 66074 86998 66076 87050
rect 66020 86996 66076 86998
rect 66124 87050 66180 87052
rect 66124 86998 66126 87050
rect 66126 86998 66178 87050
rect 66178 86998 66180 87050
rect 66124 86996 66180 86998
rect 65916 85482 65972 85484
rect 65916 85430 65918 85482
rect 65918 85430 65970 85482
rect 65970 85430 65972 85482
rect 65916 85428 65972 85430
rect 66020 85482 66076 85484
rect 66020 85430 66022 85482
rect 66022 85430 66074 85482
rect 66074 85430 66076 85482
rect 66020 85428 66076 85430
rect 66124 85482 66180 85484
rect 66124 85430 66126 85482
rect 66126 85430 66178 85482
rect 66178 85430 66180 85482
rect 66124 85428 66180 85430
rect 65916 83914 65972 83916
rect 65916 83862 65918 83914
rect 65918 83862 65970 83914
rect 65970 83862 65972 83914
rect 65916 83860 65972 83862
rect 66020 83914 66076 83916
rect 66020 83862 66022 83914
rect 66022 83862 66074 83914
rect 66074 83862 66076 83914
rect 66020 83860 66076 83862
rect 66124 83914 66180 83916
rect 66124 83862 66126 83914
rect 66126 83862 66178 83914
rect 66178 83862 66180 83914
rect 66124 83860 66180 83862
rect 65916 82346 65972 82348
rect 65916 82294 65918 82346
rect 65918 82294 65970 82346
rect 65970 82294 65972 82346
rect 65916 82292 65972 82294
rect 66020 82346 66076 82348
rect 66020 82294 66022 82346
rect 66022 82294 66074 82346
rect 66074 82294 66076 82346
rect 66020 82292 66076 82294
rect 66124 82346 66180 82348
rect 66124 82294 66126 82346
rect 66126 82294 66178 82346
rect 66178 82294 66180 82346
rect 66124 82292 66180 82294
rect 65916 80778 65972 80780
rect 65916 80726 65918 80778
rect 65918 80726 65970 80778
rect 65970 80726 65972 80778
rect 65916 80724 65972 80726
rect 66020 80778 66076 80780
rect 66020 80726 66022 80778
rect 66022 80726 66074 80778
rect 66074 80726 66076 80778
rect 66020 80724 66076 80726
rect 66124 80778 66180 80780
rect 66124 80726 66126 80778
rect 66126 80726 66178 80778
rect 66178 80726 66180 80778
rect 66124 80724 66180 80726
rect 65916 79210 65972 79212
rect 65916 79158 65918 79210
rect 65918 79158 65970 79210
rect 65970 79158 65972 79210
rect 65916 79156 65972 79158
rect 66020 79210 66076 79212
rect 66020 79158 66022 79210
rect 66022 79158 66074 79210
rect 66074 79158 66076 79210
rect 66020 79156 66076 79158
rect 66124 79210 66180 79212
rect 66124 79158 66126 79210
rect 66126 79158 66178 79210
rect 66178 79158 66180 79210
rect 66124 79156 66180 79158
rect 65916 77642 65972 77644
rect 65916 77590 65918 77642
rect 65918 77590 65970 77642
rect 65970 77590 65972 77642
rect 65916 77588 65972 77590
rect 66020 77642 66076 77644
rect 66020 77590 66022 77642
rect 66022 77590 66074 77642
rect 66074 77590 66076 77642
rect 66020 77588 66076 77590
rect 66124 77642 66180 77644
rect 66124 77590 66126 77642
rect 66126 77590 66178 77642
rect 66178 77590 66180 77642
rect 66124 77588 66180 77590
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 67340 68012 67396 68068
rect 65324 67058 65380 67060
rect 65324 67006 65326 67058
rect 65326 67006 65378 67058
rect 65378 67006 65380 67058
rect 65324 67004 65380 67006
rect 65660 67004 65716 67060
rect 65324 65996 65380 66052
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 67116 66108 67172 66164
rect 65884 65996 65940 66052
rect 66332 66050 66388 66052
rect 66332 65998 66334 66050
rect 66334 65998 66386 66050
rect 66386 65998 66388 66050
rect 66332 65996 66388 65998
rect 65660 65548 65716 65604
rect 66780 65548 66836 65604
rect 65772 65212 65828 65268
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 65996 64706 66052 64708
rect 65996 64654 65998 64706
rect 65998 64654 66050 64706
rect 66050 64654 66052 64706
rect 65996 64652 66052 64654
rect 65436 64482 65492 64484
rect 65436 64430 65438 64482
rect 65438 64430 65490 64482
rect 65490 64430 65492 64482
rect 65436 64428 65492 64430
rect 66444 64428 66500 64484
rect 65548 64316 65604 64372
rect 65660 64034 65716 64036
rect 65660 63982 65662 64034
rect 65662 63982 65714 64034
rect 65714 63982 65716 64034
rect 65660 63980 65716 63982
rect 65324 63922 65380 63924
rect 65324 63870 65326 63922
rect 65326 63870 65378 63922
rect 65378 63870 65380 63922
rect 65324 63868 65380 63870
rect 65548 63756 65604 63812
rect 66220 63810 66276 63812
rect 66220 63758 66222 63810
rect 66222 63758 66274 63810
rect 66274 63758 66276 63810
rect 66220 63756 66276 63758
rect 65548 63532 65604 63588
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66332 63532 66388 63588
rect 66124 63476 66180 63478
rect 65436 62860 65492 62916
rect 64988 60732 65044 60788
rect 63868 60060 63924 60116
rect 64092 60396 64148 60452
rect 63532 59106 63588 59108
rect 63532 59054 63534 59106
rect 63534 59054 63586 59106
rect 63586 59054 63588 59106
rect 63532 59052 63588 59054
rect 63980 59106 64036 59108
rect 63980 59054 63982 59106
rect 63982 59054 64034 59106
rect 64034 59054 64036 59106
rect 63980 59052 64036 59054
rect 64876 60620 64932 60676
rect 64428 60060 64484 60116
rect 64764 58828 64820 58884
rect 63756 58322 63812 58324
rect 63756 58270 63758 58322
rect 63758 58270 63810 58322
rect 63810 58270 63812 58322
rect 63756 58268 63812 58270
rect 63532 57036 63588 57092
rect 63980 56924 64036 56980
rect 63532 56476 63588 56532
rect 63756 56194 63812 56196
rect 63756 56142 63758 56194
rect 63758 56142 63810 56194
rect 63810 56142 63812 56194
rect 63756 56140 63812 56142
rect 63644 55356 63700 55412
rect 63756 55916 63812 55972
rect 63644 55020 63700 55076
rect 64540 57820 64596 57876
rect 64652 57484 64708 57540
rect 64316 56866 64372 56868
rect 64316 56814 64318 56866
rect 64318 56814 64370 56866
rect 64370 56814 64372 56866
rect 64316 56812 64372 56814
rect 64092 56252 64148 56308
rect 64316 56476 64372 56532
rect 63980 55468 64036 55524
rect 64204 56140 64260 56196
rect 63532 53452 63588 53508
rect 63868 54684 63924 54740
rect 63420 52332 63476 52388
rect 63196 50652 63252 50708
rect 63084 48914 63140 48916
rect 63084 48862 63086 48914
rect 63086 48862 63138 48914
rect 63138 48862 63140 48914
rect 63084 48860 63140 48862
rect 62860 48188 62916 48244
rect 63084 48636 63140 48692
rect 63084 48300 63140 48356
rect 63084 47964 63140 48020
rect 62300 46844 62356 46900
rect 61628 44380 61684 44436
rect 61740 44940 61796 44996
rect 61516 44156 61572 44212
rect 61628 44098 61684 44100
rect 61628 44046 61630 44098
rect 61630 44046 61682 44098
rect 61682 44046 61684 44098
rect 61628 44044 61684 44046
rect 62972 47682 63028 47684
rect 62972 47630 62974 47682
rect 62974 47630 63026 47682
rect 63026 47630 63028 47682
rect 62972 47628 63028 47630
rect 64540 55916 64596 55972
rect 64652 55468 64708 55524
rect 64876 58322 64932 58324
rect 64876 58270 64878 58322
rect 64878 58270 64930 58322
rect 64930 58270 64932 58322
rect 64876 58268 64932 58270
rect 64988 56924 65044 56980
rect 64428 54738 64484 54740
rect 64428 54686 64430 54738
rect 64430 54686 64482 54738
rect 64482 54686 64484 54738
rect 64428 54684 64484 54686
rect 64876 55580 64932 55636
rect 64204 53116 64260 53172
rect 63756 52780 63812 52836
rect 64428 52274 64484 52276
rect 64428 52222 64430 52274
rect 64430 52222 64482 52274
rect 64482 52222 64484 52274
rect 64428 52220 64484 52222
rect 63868 51324 63924 51380
rect 63756 50652 63812 50708
rect 63420 49868 63476 49924
rect 63420 48972 63476 49028
rect 63308 48242 63364 48244
rect 63308 48190 63310 48242
rect 63310 48190 63362 48242
rect 63362 48190 63364 48242
rect 63308 48188 63364 48190
rect 63420 48076 63476 48132
rect 63196 46786 63252 46788
rect 63196 46734 63198 46786
rect 63198 46734 63250 46786
rect 63250 46734 63252 46786
rect 63196 46732 63252 46734
rect 62972 46674 63028 46676
rect 62972 46622 62974 46674
rect 62974 46622 63026 46674
rect 63026 46622 63028 46674
rect 62972 46620 63028 46622
rect 63084 46508 63140 46564
rect 62860 45724 62916 45780
rect 62860 45388 62916 45444
rect 61964 44546 62020 44548
rect 61964 44494 61966 44546
rect 61966 44494 62018 44546
rect 62018 44494 62020 44546
rect 61964 44492 62020 44494
rect 61740 43596 61796 43652
rect 61180 43484 61236 43540
rect 60508 42924 60564 42980
rect 60620 43036 60676 43092
rect 60172 42028 60228 42084
rect 60284 41244 60340 41300
rect 59948 5964 60004 6020
rect 60060 32732 60116 32788
rect 56588 4338 56644 4340
rect 56588 4286 56590 4338
rect 56590 4286 56642 4338
rect 56642 4286 56644 4338
rect 56588 4284 56644 4286
rect 59836 4508 59892 4564
rect 57372 4284 57428 4340
rect 59500 4396 59556 4452
rect 55468 4226 55524 4228
rect 55468 4174 55470 4226
rect 55470 4174 55522 4226
rect 55522 4174 55524 4226
rect 55468 4172 55524 4174
rect 55468 3388 55524 3444
rect 55804 3442 55860 3444
rect 55804 3390 55806 3442
rect 55806 3390 55858 3442
rect 55858 3390 55860 3442
rect 55804 3388 55860 3390
rect 56588 3442 56644 3444
rect 56588 3390 56590 3442
rect 56590 3390 56642 3442
rect 56642 3390 56644 3442
rect 56588 3388 56644 3390
rect 59500 3666 59556 3668
rect 59500 3614 59502 3666
rect 59502 3614 59554 3666
rect 59554 3614 59556 3666
rect 59500 3612 59556 3614
rect 60396 32844 60452 32900
rect 60508 40236 60564 40292
rect 60172 23772 60228 23828
rect 61180 41916 61236 41972
rect 61292 43036 61348 43092
rect 61180 41244 61236 41300
rect 61180 40572 61236 40628
rect 61516 42924 61572 42980
rect 61404 42642 61460 42644
rect 61404 42590 61406 42642
rect 61406 42590 61458 42642
rect 61458 42590 61460 42642
rect 61404 42588 61460 42590
rect 61404 41298 61460 41300
rect 61404 41246 61406 41298
rect 61406 41246 61458 41298
rect 61458 41246 61460 41298
rect 61404 41244 61460 41246
rect 61964 43820 62020 43876
rect 62188 44268 62244 44324
rect 62412 44322 62468 44324
rect 62412 44270 62414 44322
rect 62414 44270 62466 44322
rect 62466 44270 62468 44322
rect 62412 44268 62468 44270
rect 62300 43708 62356 43764
rect 61852 43372 61908 43428
rect 61628 42642 61684 42644
rect 61628 42590 61630 42642
rect 61630 42590 61682 42642
rect 61682 42590 61684 42642
rect 61628 42588 61684 42590
rect 62412 43260 62468 43316
rect 61852 42028 61908 42084
rect 61628 40962 61684 40964
rect 61628 40910 61630 40962
rect 61630 40910 61682 40962
rect 61682 40910 61684 40962
rect 61628 40908 61684 40910
rect 61964 40626 62020 40628
rect 61964 40574 61966 40626
rect 61966 40574 62018 40626
rect 62018 40574 62020 40626
rect 61964 40572 62020 40574
rect 61516 40402 61572 40404
rect 61516 40350 61518 40402
rect 61518 40350 61570 40402
rect 61570 40350 61572 40402
rect 61516 40348 61572 40350
rect 62412 40402 62468 40404
rect 62412 40350 62414 40402
rect 62414 40350 62466 40402
rect 62466 40350 62468 40402
rect 62412 40348 62468 40350
rect 62748 44492 62804 44548
rect 62748 43538 62804 43540
rect 62748 43486 62750 43538
rect 62750 43486 62802 43538
rect 62802 43486 62804 43538
rect 62748 43484 62804 43486
rect 64540 52108 64596 52164
rect 66556 64316 66612 64372
rect 66668 63756 66724 63812
rect 68908 69132 68964 69188
rect 70140 115388 70196 115444
rect 72044 116284 72100 116340
rect 71708 115666 71764 115668
rect 71708 115614 71710 115666
rect 71710 115614 71762 115666
rect 71762 115614 71764 115666
rect 71708 115612 71764 115614
rect 67340 64764 67396 64820
rect 68012 64818 68068 64820
rect 68012 64766 68014 64818
rect 68014 64766 68066 64818
rect 68066 64766 68068 64818
rect 68012 64764 68068 64766
rect 67116 63980 67172 64036
rect 67340 64428 67396 64484
rect 66780 63196 66836 63252
rect 65772 62860 65828 62916
rect 68124 64428 68180 64484
rect 67564 63868 67620 63924
rect 67452 63810 67508 63812
rect 67452 63758 67454 63810
rect 67454 63758 67506 63810
rect 67506 63758 67508 63810
rect 67452 63756 67508 63758
rect 67340 62524 67396 62580
rect 67676 64092 67732 64148
rect 68012 63250 68068 63252
rect 68012 63198 68014 63250
rect 68014 63198 68066 63250
rect 68066 63198 68068 63250
rect 68012 63196 68068 63198
rect 67564 62412 67620 62468
rect 65660 62354 65716 62356
rect 65660 62302 65662 62354
rect 65662 62302 65714 62354
rect 65714 62302 65716 62354
rect 65660 62300 65716 62302
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65212 60620 65268 60676
rect 65324 60732 65380 60788
rect 65436 60562 65492 60564
rect 65436 60510 65438 60562
rect 65438 60510 65490 60562
rect 65490 60510 65492 60562
rect 65436 60508 65492 60510
rect 65660 60508 65716 60564
rect 65324 58828 65380 58884
rect 65548 59052 65604 59108
rect 65548 58268 65604 58324
rect 65436 57484 65492 57540
rect 65324 57090 65380 57092
rect 65324 57038 65326 57090
rect 65326 57038 65378 57090
rect 65378 57038 65380 57090
rect 65324 57036 65380 57038
rect 65548 57148 65604 57204
rect 65548 56978 65604 56980
rect 65548 56926 65550 56978
rect 65550 56926 65602 56978
rect 65602 56926 65604 56978
rect 65548 56924 65604 56926
rect 65548 56476 65604 56532
rect 65548 55580 65604 55636
rect 65100 55132 65156 55188
rect 65100 54236 65156 54292
rect 65436 53676 65492 53732
rect 66332 61292 66388 61348
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65884 59106 65940 59108
rect 65884 59054 65886 59106
rect 65886 59054 65938 59106
rect 65938 59054 65940 59106
rect 65884 59052 65940 59054
rect 67452 61852 67508 61908
rect 66668 61570 66724 61572
rect 66668 61518 66670 61570
rect 66670 61518 66722 61570
rect 66722 61518 66724 61570
rect 66668 61516 66724 61518
rect 67228 61516 67284 61572
rect 66668 60674 66724 60676
rect 66668 60622 66670 60674
rect 66670 60622 66722 60674
rect 66722 60622 66724 60674
rect 66668 60620 66724 60622
rect 67900 61628 67956 61684
rect 67340 61346 67396 61348
rect 67340 61294 67342 61346
rect 67342 61294 67394 61346
rect 67394 61294 67396 61346
rect 67340 61292 67396 61294
rect 67676 61068 67732 61124
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65772 58322 65828 58324
rect 65772 58270 65774 58322
rect 65774 58270 65826 58322
rect 65826 58270 65828 58322
rect 65772 58268 65828 58270
rect 65884 58156 65940 58212
rect 66220 58210 66276 58212
rect 66220 58158 66222 58210
rect 66222 58158 66274 58210
rect 66274 58158 66276 58210
rect 66220 58156 66276 58158
rect 65772 57650 65828 57652
rect 65772 57598 65774 57650
rect 65774 57598 65826 57650
rect 65826 57598 65828 57650
rect 65772 57596 65828 57598
rect 66332 57596 66388 57652
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 66780 60284 66836 60340
rect 66780 59164 66836 59220
rect 66556 57596 66612 57652
rect 66668 59052 66724 59108
rect 66444 56924 66500 56980
rect 66668 57036 66724 57092
rect 67228 60508 67284 60564
rect 67004 60396 67060 60452
rect 67564 60620 67620 60676
rect 68124 61068 68180 61124
rect 68012 60898 68068 60900
rect 68012 60846 68014 60898
rect 68014 60846 68066 60898
rect 68066 60846 68068 60898
rect 68012 60844 68068 60846
rect 67900 60396 67956 60452
rect 67116 59106 67172 59108
rect 67116 59054 67118 59106
rect 67118 59054 67170 59106
rect 67170 59054 67172 59106
rect 67116 59052 67172 59054
rect 67004 58828 67060 58884
rect 67676 58940 67732 58996
rect 67228 58434 67284 58436
rect 67228 58382 67230 58434
rect 67230 58382 67282 58434
rect 67282 58382 67284 58434
rect 67228 58380 67284 58382
rect 66892 56812 66948 56868
rect 66332 56588 66388 56644
rect 65772 55970 65828 55972
rect 65772 55918 65774 55970
rect 65774 55918 65826 55970
rect 65826 55918 65828 55970
rect 65772 55916 65828 55918
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65996 55410 66052 55412
rect 65996 55358 65998 55410
rect 65998 55358 66050 55410
rect 66050 55358 66052 55410
rect 65996 55356 66052 55358
rect 67004 56700 67060 56756
rect 66668 56588 66724 56644
rect 66556 55692 66612 55748
rect 66668 55356 66724 55412
rect 66332 54684 66388 54740
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65660 53564 65716 53620
rect 64988 52332 65044 52388
rect 64988 52050 65044 52052
rect 64988 51998 64990 52050
rect 64990 51998 65042 52050
rect 65042 51998 65044 52050
rect 64988 51996 65044 51998
rect 63980 51100 64036 51156
rect 63980 50764 64036 50820
rect 64876 51660 64932 51716
rect 64540 50988 64596 51044
rect 64316 50482 64372 50484
rect 64316 50430 64318 50482
rect 64318 50430 64370 50482
rect 64370 50430 64372 50482
rect 64316 50428 64372 50430
rect 64204 49922 64260 49924
rect 64204 49870 64206 49922
rect 64206 49870 64258 49922
rect 64258 49870 64260 49922
rect 64204 49868 64260 49870
rect 64876 50988 64932 51044
rect 65436 52050 65492 52052
rect 65436 51998 65438 52050
rect 65438 51998 65490 52050
rect 65490 51998 65492 52050
rect 65436 51996 65492 51998
rect 65212 51660 65268 51716
rect 65100 51100 65156 51156
rect 65212 51324 65268 51380
rect 64988 50540 65044 50596
rect 65100 50764 65156 50820
rect 64764 50370 64820 50372
rect 64764 50318 64766 50370
rect 64766 50318 64818 50370
rect 64818 50318 64820 50370
rect 64764 50316 64820 50318
rect 63980 49084 64036 49140
rect 64204 48466 64260 48468
rect 64204 48414 64206 48466
rect 64206 48414 64258 48466
rect 64258 48414 64260 48466
rect 64204 48412 64260 48414
rect 63980 48242 64036 48244
rect 63980 48190 63982 48242
rect 63982 48190 64034 48242
rect 64034 48190 64036 48242
rect 63980 48188 64036 48190
rect 64316 48076 64372 48132
rect 64204 47628 64260 47684
rect 63532 46732 63588 46788
rect 63980 47516 64036 47572
rect 63756 46674 63812 46676
rect 63756 46622 63758 46674
rect 63758 46622 63810 46674
rect 63810 46622 63812 46674
rect 63756 46620 63812 46622
rect 63868 45778 63924 45780
rect 63868 45726 63870 45778
rect 63870 45726 63922 45778
rect 63922 45726 63924 45778
rect 63868 45724 63924 45726
rect 63532 45276 63588 45332
rect 63308 44492 63364 44548
rect 62972 44210 63028 44212
rect 62972 44158 62974 44210
rect 62974 44158 63026 44210
rect 63026 44158 63028 44210
rect 62972 44156 63028 44158
rect 63420 44156 63476 44212
rect 63196 44044 63252 44100
rect 63084 43650 63140 43652
rect 63084 43598 63086 43650
rect 63086 43598 63138 43650
rect 63138 43598 63140 43650
rect 63084 43596 63140 43598
rect 63084 43372 63140 43428
rect 64092 47292 64148 47348
rect 64092 45836 64148 45892
rect 64316 46956 64372 47012
rect 64540 48412 64596 48468
rect 64316 45164 64372 45220
rect 64540 45330 64596 45332
rect 64540 45278 64542 45330
rect 64542 45278 64594 45330
rect 64594 45278 64596 45330
rect 64540 45276 64596 45278
rect 65436 50652 65492 50708
rect 66332 53900 66388 53956
rect 66220 53340 66276 53396
rect 66556 54626 66612 54628
rect 66556 54574 66558 54626
rect 66558 54574 66610 54626
rect 66610 54574 66612 54626
rect 66556 54572 66612 54574
rect 67004 54572 67060 54628
rect 66556 54012 66612 54068
rect 66892 54460 66948 54516
rect 67004 53954 67060 53956
rect 67004 53902 67006 53954
rect 67006 53902 67058 53954
rect 67058 53902 67060 53954
rect 67004 53900 67060 53902
rect 66444 53452 66500 53508
rect 67004 53228 67060 53284
rect 66332 52946 66388 52948
rect 66332 52894 66334 52946
rect 66334 52894 66386 52946
rect 66386 52894 66388 52946
rect 66332 52892 66388 52894
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65884 52332 65940 52388
rect 66668 52332 66724 52388
rect 66220 51660 66276 51716
rect 65884 51324 65940 51380
rect 65660 50594 65716 50596
rect 65660 50542 65662 50594
rect 65662 50542 65714 50594
rect 65714 50542 65716 50594
rect 65660 50540 65716 50542
rect 65324 50316 65380 50372
rect 65324 49698 65380 49700
rect 65324 49646 65326 49698
rect 65326 49646 65378 49698
rect 65378 49646 65380 49698
rect 65324 49644 65380 49646
rect 65324 48636 65380 48692
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65772 49196 65828 49252
rect 63980 44156 64036 44212
rect 64204 44210 64260 44212
rect 64204 44158 64206 44210
rect 64206 44158 64258 44210
rect 64258 44158 64260 44210
rect 64204 44156 64260 44158
rect 63532 43708 63588 43764
rect 63868 43820 63924 43876
rect 63532 42642 63588 42644
rect 63532 42590 63534 42642
rect 63534 42590 63586 42642
rect 63586 42590 63588 42642
rect 63532 42588 63588 42590
rect 64204 43820 64260 43876
rect 64540 43820 64596 43876
rect 63980 42812 64036 42868
rect 64428 43260 64484 43316
rect 65548 48076 65604 48132
rect 65324 44492 65380 44548
rect 65324 43538 65380 43540
rect 65324 43486 65326 43538
rect 65326 43486 65378 43538
rect 65378 43486 65380 43538
rect 65324 43484 65380 43486
rect 65212 43260 65268 43316
rect 63980 42028 64036 42084
rect 62748 40962 62804 40964
rect 62748 40910 62750 40962
rect 62750 40910 62802 40962
rect 62802 40910 62804 40962
rect 62748 40908 62804 40910
rect 65772 48018 65828 48020
rect 65772 47966 65774 48018
rect 65774 47966 65826 48018
rect 65826 47966 65828 48018
rect 65772 47964 65828 47966
rect 66108 47964 66164 48020
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 66556 51548 66612 51604
rect 67452 56642 67508 56644
rect 67452 56590 67454 56642
rect 67454 56590 67506 56642
rect 67506 56590 67508 56642
rect 67452 56588 67508 56590
rect 67340 55692 67396 55748
rect 67452 54348 67508 54404
rect 67340 54012 67396 54068
rect 67452 53676 67508 53732
rect 66780 51996 66836 52052
rect 67004 51548 67060 51604
rect 67228 51772 67284 51828
rect 67116 50764 67172 50820
rect 67452 52220 67508 52276
rect 67900 56866 67956 56868
rect 67900 56814 67902 56866
rect 67902 56814 67954 56866
rect 67954 56814 67956 56866
rect 67900 56812 67956 56814
rect 67788 56476 67844 56532
rect 67788 55804 67844 55860
rect 68460 64706 68516 64708
rect 68460 64654 68462 64706
rect 68462 64654 68514 64706
rect 68514 64654 68516 64706
rect 68460 64652 68516 64654
rect 68572 64092 68628 64148
rect 69020 63532 69076 63588
rect 69356 64706 69412 64708
rect 69356 64654 69358 64706
rect 69358 64654 69410 64706
rect 69410 64654 69412 64706
rect 69356 64652 69412 64654
rect 70252 66780 70308 66836
rect 70700 66444 70756 66500
rect 70476 65996 70532 66052
rect 70476 64876 70532 64932
rect 70700 65548 70756 65604
rect 69132 63196 69188 63252
rect 69916 64594 69972 64596
rect 69916 64542 69918 64594
rect 69918 64542 69970 64594
rect 69970 64542 69972 64594
rect 69916 64540 69972 64542
rect 70588 64594 70644 64596
rect 70588 64542 70590 64594
rect 70590 64542 70642 64594
rect 70642 64542 70644 64594
rect 70588 64540 70644 64542
rect 70476 64428 70532 64484
rect 70700 64146 70756 64148
rect 70700 64094 70702 64146
rect 70702 64094 70754 64146
rect 70754 64094 70756 64146
rect 70700 64092 70756 64094
rect 69468 63922 69524 63924
rect 69468 63870 69470 63922
rect 69470 63870 69522 63922
rect 69522 63870 69524 63922
rect 69468 63868 69524 63870
rect 70476 63922 70532 63924
rect 70476 63870 70478 63922
rect 70478 63870 70530 63922
rect 70530 63870 70532 63922
rect 70476 63868 70532 63870
rect 70140 63420 70196 63476
rect 68572 62972 68628 63028
rect 68460 62914 68516 62916
rect 68460 62862 68462 62914
rect 68462 62862 68514 62914
rect 68514 62862 68516 62914
rect 68460 62860 68516 62862
rect 69356 63026 69412 63028
rect 69356 62974 69358 63026
rect 69358 62974 69410 63026
rect 69410 62974 69412 63026
rect 69356 62972 69412 62974
rect 69468 62914 69524 62916
rect 69468 62862 69470 62914
rect 69470 62862 69522 62914
rect 69522 62862 69524 62914
rect 69468 62860 69524 62862
rect 70140 62972 70196 63028
rect 69580 62242 69636 62244
rect 69580 62190 69582 62242
rect 69582 62190 69634 62242
rect 69634 62190 69636 62242
rect 69580 62188 69636 62190
rect 68348 61682 68404 61684
rect 68348 61630 68350 61682
rect 68350 61630 68402 61682
rect 68402 61630 68404 61682
rect 68348 61628 68404 61630
rect 68572 61010 68628 61012
rect 68572 60958 68574 61010
rect 68574 60958 68626 61010
rect 68626 60958 68628 61010
rect 68572 60956 68628 60958
rect 68684 60396 68740 60452
rect 68572 59500 68628 59556
rect 68348 59388 68404 59444
rect 68460 59106 68516 59108
rect 68460 59054 68462 59106
rect 68462 59054 68514 59106
rect 68514 59054 68516 59106
rect 68460 59052 68516 59054
rect 68572 58940 68628 58996
rect 68460 58828 68516 58884
rect 68572 58546 68628 58548
rect 68572 58494 68574 58546
rect 68574 58494 68626 58546
rect 68626 58494 68628 58546
rect 68572 58492 68628 58494
rect 70028 62578 70084 62580
rect 70028 62526 70030 62578
rect 70030 62526 70082 62578
rect 70082 62526 70084 62578
rect 70028 62524 70084 62526
rect 70028 61852 70084 61908
rect 70364 61628 70420 61684
rect 70028 61346 70084 61348
rect 70028 61294 70030 61346
rect 70030 61294 70082 61346
rect 70082 61294 70084 61346
rect 70028 61292 70084 61294
rect 69356 60956 69412 61012
rect 69804 60786 69860 60788
rect 69804 60734 69806 60786
rect 69806 60734 69858 60786
rect 69858 60734 69860 60786
rect 69804 60732 69860 60734
rect 69468 60508 69524 60564
rect 69356 60172 69412 60228
rect 70252 60844 70308 60900
rect 70476 60956 70532 61012
rect 70364 60172 70420 60228
rect 69580 59948 69636 60004
rect 68908 59500 68964 59556
rect 69356 59442 69412 59444
rect 69356 59390 69358 59442
rect 69358 59390 69410 59442
rect 69410 59390 69412 59442
rect 69356 59388 69412 59390
rect 69468 59218 69524 59220
rect 69468 59166 69470 59218
rect 69470 59166 69522 59218
rect 69522 59166 69524 59218
rect 69468 59164 69524 59166
rect 69356 59052 69412 59108
rect 69132 58828 69188 58884
rect 69692 59500 69748 59556
rect 69580 58940 69636 58996
rect 70028 59724 70084 59780
rect 69916 59442 69972 59444
rect 69916 59390 69918 59442
rect 69918 59390 69970 59442
rect 69970 59390 69972 59442
rect 69916 59388 69972 59390
rect 70028 59052 70084 59108
rect 69804 58604 69860 58660
rect 69916 58940 69972 58996
rect 69580 58492 69636 58548
rect 69244 58380 69300 58436
rect 69468 58380 69524 58436
rect 68572 56476 68628 56532
rect 68572 56306 68628 56308
rect 68572 56254 68574 56306
rect 68574 56254 68626 56306
rect 68626 56254 68628 56306
rect 68572 56252 68628 56254
rect 70028 58828 70084 58884
rect 70588 62188 70644 62244
rect 72380 115666 72436 115668
rect 72380 115614 72382 115666
rect 72382 115614 72434 115666
rect 72434 115614 72436 115666
rect 72380 115612 72436 115614
rect 71260 94386 71316 94388
rect 71260 94334 71262 94386
rect 71262 94334 71314 94386
rect 71314 94334 71316 94386
rect 71260 94332 71316 94334
rect 71820 94386 71876 94388
rect 71820 94334 71822 94386
rect 71822 94334 71874 94386
rect 71874 94334 71876 94386
rect 71820 94332 71876 94334
rect 72156 94274 72212 94276
rect 72156 94222 72158 94274
rect 72158 94222 72210 94274
rect 72210 94222 72212 94274
rect 72156 94220 72212 94222
rect 72380 68124 72436 68180
rect 71708 66444 71764 66500
rect 71260 64482 71316 64484
rect 71260 64430 71262 64482
rect 71262 64430 71314 64482
rect 71314 64430 71316 64482
rect 71260 64428 71316 64430
rect 71148 64092 71204 64148
rect 71148 63922 71204 63924
rect 71148 63870 71150 63922
rect 71150 63870 71202 63922
rect 71202 63870 71204 63922
rect 71148 63868 71204 63870
rect 71148 62300 71204 62356
rect 70924 62242 70980 62244
rect 70924 62190 70926 62242
rect 70926 62190 70978 62242
rect 70978 62190 70980 62242
rect 70924 62188 70980 62190
rect 70812 61852 70868 61908
rect 71148 61628 71204 61684
rect 70588 59388 70644 59444
rect 70700 61292 70756 61348
rect 70364 58828 70420 58884
rect 70924 60898 70980 60900
rect 70924 60846 70926 60898
rect 70926 60846 70978 60898
rect 70978 60846 70980 60898
rect 70924 60844 70980 60846
rect 71372 62300 71428 62356
rect 71484 64428 71540 64484
rect 71708 64482 71764 64484
rect 71708 64430 71710 64482
rect 71710 64430 71762 64482
rect 71762 64430 71764 64482
rect 71708 64428 71764 64430
rect 71708 62354 71764 62356
rect 71708 62302 71710 62354
rect 71710 62302 71762 62354
rect 71762 62302 71764 62354
rect 71708 62300 71764 62302
rect 71708 61292 71764 61348
rect 70924 59778 70980 59780
rect 70924 59726 70926 59778
rect 70926 59726 70978 59778
rect 70978 59726 70980 59778
rect 70924 59724 70980 59726
rect 70812 59164 70868 59220
rect 71148 59724 71204 59780
rect 70924 58380 70980 58436
rect 69580 56924 69636 56980
rect 69132 56476 69188 56532
rect 68460 55916 68516 55972
rect 68348 55804 68404 55860
rect 68124 55356 68180 55412
rect 68012 54796 68068 54852
rect 72156 67116 72212 67172
rect 72380 67172 72436 67228
rect 72268 67004 72324 67060
rect 72380 66780 72436 66836
rect 72156 65548 72212 65604
rect 72380 62354 72436 62356
rect 72380 62302 72382 62354
rect 72382 62302 72434 62354
rect 72434 62302 72436 62354
rect 72380 62300 72436 62302
rect 72044 61628 72100 61684
rect 72156 61852 72212 61908
rect 71932 61010 71988 61012
rect 71932 60958 71934 61010
rect 71934 60958 71986 61010
rect 71986 60958 71988 61010
rect 71932 60956 71988 60958
rect 71932 60786 71988 60788
rect 71932 60734 71934 60786
rect 71934 60734 71986 60786
rect 71986 60734 71988 60786
rect 71932 60732 71988 60734
rect 71260 58210 71316 58212
rect 71260 58158 71262 58210
rect 71262 58158 71314 58210
rect 71314 58158 71316 58210
rect 71260 58156 71316 58158
rect 71372 58044 71428 58100
rect 71484 59500 71540 59556
rect 69692 56252 69748 56308
rect 70140 56252 70196 56308
rect 68908 56082 68964 56084
rect 68908 56030 68910 56082
rect 68910 56030 68962 56082
rect 68962 56030 68964 56082
rect 68908 56028 68964 56030
rect 68460 54796 68516 54852
rect 69356 55468 69412 55524
rect 68684 55132 68740 55188
rect 68124 54348 68180 54404
rect 68236 53506 68292 53508
rect 68236 53454 68238 53506
rect 68238 53454 68290 53506
rect 68290 53454 68292 53506
rect 68236 53452 68292 53454
rect 68012 53116 68068 53172
rect 68908 55244 68964 55300
rect 68796 54572 68852 54628
rect 67676 52108 67732 52164
rect 67228 50706 67284 50708
rect 67228 50654 67230 50706
rect 67230 50654 67282 50706
rect 67282 50654 67284 50706
rect 67228 50652 67284 50654
rect 66444 49756 66500 49812
rect 66780 49644 66836 49700
rect 66444 48748 66500 48804
rect 66780 49196 66836 49252
rect 66332 47628 66388 47684
rect 66220 47346 66276 47348
rect 66220 47294 66222 47346
rect 66222 47294 66274 47346
rect 66274 47294 66276 47346
rect 66220 47292 66276 47294
rect 66668 48130 66724 48132
rect 66668 48078 66670 48130
rect 66670 48078 66722 48130
rect 66722 48078 66724 48130
rect 66668 48076 66724 48078
rect 66668 47516 66724 47572
rect 66444 47292 66500 47348
rect 66668 46956 66724 47012
rect 65772 46898 65828 46900
rect 65772 46846 65774 46898
rect 65774 46846 65826 46898
rect 65826 46846 65828 46898
rect 65772 46844 65828 46846
rect 66220 46786 66276 46788
rect 66220 46734 66222 46786
rect 66222 46734 66274 46786
rect 66274 46734 66276 46786
rect 66220 46732 66276 46734
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65772 45218 65828 45220
rect 65772 45166 65774 45218
rect 65774 45166 65826 45218
rect 65826 45166 65828 45218
rect 65772 45164 65828 45166
rect 66444 44828 66500 44884
rect 66892 48636 66948 48692
rect 67116 48300 67172 48356
rect 67564 51602 67620 51604
rect 67564 51550 67566 51602
rect 67566 51550 67618 51602
rect 67618 51550 67620 51602
rect 67564 51548 67620 51550
rect 67788 50594 67844 50596
rect 67788 50542 67790 50594
rect 67790 50542 67842 50594
rect 67842 50542 67844 50594
rect 67788 50540 67844 50542
rect 67676 50316 67732 50372
rect 68012 51436 68068 51492
rect 68124 51378 68180 51380
rect 68124 51326 68126 51378
rect 68126 51326 68178 51378
rect 68178 51326 68180 51378
rect 68124 51324 68180 51326
rect 68124 49810 68180 49812
rect 68124 49758 68126 49810
rect 68126 49758 68178 49810
rect 68178 49758 68180 49810
rect 68124 49756 68180 49758
rect 68460 52220 68516 52276
rect 69692 55356 69748 55412
rect 69580 55186 69636 55188
rect 69580 55134 69582 55186
rect 69582 55134 69634 55186
rect 69634 55134 69636 55186
rect 69580 55132 69636 55134
rect 69468 55074 69524 55076
rect 69468 55022 69470 55074
rect 69470 55022 69522 55074
rect 69522 55022 69524 55074
rect 69468 55020 69524 55022
rect 68908 53788 68964 53844
rect 69132 54402 69188 54404
rect 69132 54350 69134 54402
rect 69134 54350 69186 54402
rect 69186 54350 69188 54402
rect 69132 54348 69188 54350
rect 69244 53116 69300 53172
rect 69244 52162 69300 52164
rect 69244 52110 69246 52162
rect 69246 52110 69298 52162
rect 69298 52110 69300 52162
rect 69244 52108 69300 52110
rect 68572 51772 68628 51828
rect 68572 51548 68628 51604
rect 69468 51490 69524 51492
rect 69468 51438 69470 51490
rect 69470 51438 69522 51490
rect 69522 51438 69524 51490
rect 69468 51436 69524 51438
rect 68908 51378 68964 51380
rect 68908 51326 68910 51378
rect 68910 51326 68962 51378
rect 68962 51326 68964 51378
rect 68908 51324 68964 51326
rect 68684 50764 68740 50820
rect 68572 50092 68628 50148
rect 68572 49698 68628 49700
rect 68572 49646 68574 49698
rect 68574 49646 68626 49698
rect 68626 49646 68628 49698
rect 68572 49644 68628 49646
rect 68348 49532 68404 49588
rect 67452 48972 67508 49028
rect 67452 48802 67508 48804
rect 67452 48750 67454 48802
rect 67454 48750 67506 48802
rect 67506 48750 67508 48802
rect 67452 48748 67508 48750
rect 67788 48748 67844 48804
rect 67004 47964 67060 48020
rect 67228 46562 67284 46564
rect 67228 46510 67230 46562
rect 67230 46510 67282 46562
rect 67282 46510 67284 46562
rect 67228 46508 67284 46510
rect 67452 48524 67508 48580
rect 67900 48076 67956 48132
rect 67676 47964 67732 48020
rect 67564 47346 67620 47348
rect 67564 47294 67566 47346
rect 67566 47294 67618 47346
rect 67618 47294 67620 47346
rect 67564 47292 67620 47294
rect 67788 47234 67844 47236
rect 67788 47182 67790 47234
rect 67790 47182 67842 47234
rect 67842 47182 67844 47234
rect 67788 47180 67844 47182
rect 67452 46060 67508 46116
rect 68012 46674 68068 46676
rect 68012 46622 68014 46674
rect 68014 46622 68066 46674
rect 68066 46622 68068 46674
rect 68012 46620 68068 46622
rect 68012 45778 68068 45780
rect 68012 45726 68014 45778
rect 68014 45726 68066 45778
rect 68066 45726 68068 45778
rect 68012 45724 68068 45726
rect 67004 45612 67060 45668
rect 67564 45666 67620 45668
rect 67564 45614 67566 45666
rect 67566 45614 67618 45666
rect 67618 45614 67620 45666
rect 67564 45612 67620 45614
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 66332 44604 66388 44660
rect 65660 44322 65716 44324
rect 65660 44270 65662 44322
rect 65662 44270 65714 44322
rect 65714 44270 65716 44322
rect 65660 44268 65716 44270
rect 66108 44322 66164 44324
rect 66108 44270 66110 44322
rect 66110 44270 66162 44322
rect 66162 44270 66164 44322
rect 66108 44268 66164 44270
rect 65660 43708 65716 43764
rect 66332 43820 66388 43876
rect 66668 44492 66724 44548
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65548 39788 65604 39844
rect 62636 39340 62692 39396
rect 62972 39564 63028 39620
rect 62860 38946 62916 38948
rect 62860 38894 62862 38946
rect 62862 38894 62914 38946
rect 62914 38894 62916 38946
rect 62860 38892 62916 38894
rect 60620 31948 60676 32004
rect 62748 26460 62804 26516
rect 62748 5068 62804 5124
rect 61068 4508 61124 4564
rect 60508 3612 60564 3668
rect 63420 39340 63476 39396
rect 63868 38946 63924 38948
rect 63868 38894 63870 38946
rect 63870 38894 63922 38946
rect 63922 38894 63924 38946
rect 63868 38892 63924 38894
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 67228 44828 67284 44884
rect 66892 44322 66948 44324
rect 66892 44270 66894 44322
rect 66894 44270 66946 44322
rect 66946 44270 66948 44322
rect 66892 44268 66948 44270
rect 67004 44098 67060 44100
rect 67004 44046 67006 44098
rect 67006 44046 67058 44098
rect 67058 44046 67060 44098
rect 67004 44044 67060 44046
rect 67116 43932 67172 43988
rect 67452 43708 67508 43764
rect 66780 42812 66836 42868
rect 63196 26514 63252 26516
rect 63196 26462 63198 26514
rect 63198 26462 63250 26514
rect 63250 26462 63252 26514
rect 63196 26460 63252 26462
rect 63868 23772 63924 23828
rect 64764 8034 64820 8036
rect 64764 7982 64766 8034
rect 64766 7982 64818 8034
rect 64818 7982 64820 8034
rect 64764 7980 64820 7982
rect 63980 5122 64036 5124
rect 63980 5070 63982 5122
rect 63982 5070 64034 5122
rect 64034 5070 64036 5122
rect 63980 5068 64036 5070
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 63868 3724 63924 3780
rect 63308 3388 63364 3444
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 68348 48748 68404 48804
rect 68460 48354 68516 48356
rect 68460 48302 68462 48354
rect 68462 48302 68514 48354
rect 68514 48302 68516 48354
rect 68460 48300 68516 48302
rect 68796 48242 68852 48244
rect 68796 48190 68798 48242
rect 68798 48190 68850 48242
rect 68850 48190 68852 48242
rect 68796 48188 68852 48190
rect 68348 47570 68404 47572
rect 68348 47518 68350 47570
rect 68350 47518 68402 47570
rect 68402 47518 68404 47570
rect 68348 47516 68404 47518
rect 70588 57036 70644 57092
rect 70364 55298 70420 55300
rect 70364 55246 70366 55298
rect 70366 55246 70418 55298
rect 70418 55246 70420 55298
rect 70364 55244 70420 55246
rect 69692 54348 69748 54404
rect 70140 54236 70196 54292
rect 70028 53730 70084 53732
rect 70028 53678 70030 53730
rect 70030 53678 70082 53730
rect 70082 53678 70084 53730
rect 70028 53676 70084 53678
rect 69692 52780 69748 52836
rect 69692 52332 69748 52388
rect 70700 56252 70756 56308
rect 70588 55298 70644 55300
rect 70588 55246 70590 55298
rect 70590 55246 70642 55298
rect 70642 55246 70644 55298
rect 70588 55244 70644 55246
rect 70476 54402 70532 54404
rect 70476 54350 70478 54402
rect 70478 54350 70530 54402
rect 70530 54350 70532 54402
rect 70476 54348 70532 54350
rect 70252 52220 70308 52276
rect 69916 51324 69972 51380
rect 69916 50428 69972 50484
rect 70588 53004 70644 53060
rect 70476 51266 70532 51268
rect 70476 51214 70478 51266
rect 70478 51214 70530 51266
rect 70530 51214 70532 51266
rect 70476 51212 70532 51214
rect 70700 52834 70756 52836
rect 70700 52782 70702 52834
rect 70702 52782 70754 52834
rect 70754 52782 70756 52834
rect 70700 52780 70756 52782
rect 70700 52220 70756 52276
rect 70924 56978 70980 56980
rect 70924 56926 70926 56978
rect 70926 56926 70978 56978
rect 70978 56926 70980 56978
rect 70924 56924 70980 56926
rect 71260 57036 71316 57092
rect 71708 58210 71764 58212
rect 71708 58158 71710 58210
rect 71710 58158 71762 58210
rect 71762 58158 71764 58210
rect 71708 58156 71764 58158
rect 71148 56252 71204 56308
rect 71036 55970 71092 55972
rect 71036 55918 71038 55970
rect 71038 55918 71090 55970
rect 71090 55918 71092 55970
rect 71036 55916 71092 55918
rect 71036 55186 71092 55188
rect 71036 55134 71038 55186
rect 71038 55134 71090 55186
rect 71090 55134 71092 55186
rect 71036 55132 71092 55134
rect 71260 53730 71316 53732
rect 71260 53678 71262 53730
rect 71262 53678 71314 53730
rect 71314 53678 71316 53730
rect 71260 53676 71316 53678
rect 70924 53506 70980 53508
rect 70924 53454 70926 53506
rect 70926 53454 70978 53506
rect 70978 53454 70980 53506
rect 70924 53452 70980 53454
rect 71596 57036 71652 57092
rect 71484 56028 71540 56084
rect 71484 55468 71540 55524
rect 71708 55356 71764 55412
rect 71484 55298 71540 55300
rect 71484 55246 71486 55298
rect 71486 55246 71538 55298
rect 71538 55246 71540 55298
rect 71484 55244 71540 55246
rect 71484 51378 71540 51380
rect 71484 51326 71486 51378
rect 71486 51326 71538 51378
rect 71538 51326 71540 51378
rect 71484 51324 71540 51326
rect 71148 51212 71204 51268
rect 72044 59442 72100 59444
rect 72044 59390 72046 59442
rect 72046 59390 72098 59442
rect 72098 59390 72100 59442
rect 72044 59388 72100 59390
rect 72044 58044 72100 58100
rect 71932 56252 71988 56308
rect 71932 55970 71988 55972
rect 71932 55918 71934 55970
rect 71934 55918 71986 55970
rect 71986 55918 71988 55970
rect 71932 55916 71988 55918
rect 71932 55074 71988 55076
rect 71932 55022 71934 55074
rect 71934 55022 71986 55074
rect 71986 55022 71988 55074
rect 71932 55020 71988 55022
rect 72380 60956 72436 61012
rect 72268 60620 72324 60676
rect 75404 116508 75460 116564
rect 74396 116338 74452 116340
rect 74396 116286 74398 116338
rect 74398 116286 74450 116338
rect 74450 116286 74452 116338
rect 74396 116284 74452 116286
rect 75516 116226 75572 116228
rect 75516 116174 75518 116226
rect 75518 116174 75570 116226
rect 75570 116174 75572 116226
rect 75516 116172 75572 116174
rect 76188 116172 76244 116228
rect 73388 115836 73444 115892
rect 74172 115836 74228 115892
rect 74732 113372 74788 113428
rect 73948 106204 74004 106260
rect 73948 102956 74004 103012
rect 74732 93436 74788 93492
rect 74732 87276 74788 87332
rect 73276 67004 73332 67060
rect 74284 66892 74340 66948
rect 74620 66780 74676 66836
rect 73276 66444 73332 66500
rect 74172 66444 74228 66500
rect 74620 66220 74676 66276
rect 76972 116562 77028 116564
rect 76972 116510 76974 116562
rect 76974 116510 77026 116562
rect 77026 116510 77028 116562
rect 76972 116508 77028 116510
rect 78092 116508 78148 116564
rect 76748 115724 76804 115780
rect 77532 115724 77588 115780
rect 74956 66892 75012 66948
rect 74732 65884 74788 65940
rect 74172 65378 74228 65380
rect 74172 65326 74174 65378
rect 74174 65326 74226 65378
rect 74226 65326 74228 65378
rect 74172 65324 74228 65326
rect 74172 64316 74228 64372
rect 73948 64204 74004 64260
rect 73388 63644 73444 63700
rect 73388 62466 73444 62468
rect 73388 62414 73390 62466
rect 73390 62414 73442 62466
rect 73442 62414 73444 62466
rect 73388 62412 73444 62414
rect 73500 62354 73556 62356
rect 73500 62302 73502 62354
rect 73502 62302 73554 62354
rect 73554 62302 73556 62354
rect 73500 62300 73556 62302
rect 73724 62354 73780 62356
rect 73724 62302 73726 62354
rect 73726 62302 73778 62354
rect 73778 62302 73780 62354
rect 73724 62300 73780 62302
rect 73052 59778 73108 59780
rect 73052 59726 73054 59778
rect 73054 59726 73106 59778
rect 73106 59726 73108 59778
rect 73052 59724 73108 59726
rect 73500 61292 73556 61348
rect 73052 57036 73108 57092
rect 72492 56812 72548 56868
rect 73612 61010 73668 61012
rect 73612 60958 73614 61010
rect 73614 60958 73666 61010
rect 73666 60958 73668 61010
rect 73612 60956 73668 60958
rect 73612 60674 73668 60676
rect 73612 60622 73614 60674
rect 73614 60622 73666 60674
rect 73666 60622 73668 60674
rect 73612 60620 73668 60622
rect 72604 55916 72660 55972
rect 72604 54402 72660 54404
rect 72604 54350 72606 54402
rect 72606 54350 72658 54402
rect 72658 54350 72660 54402
rect 72604 54348 72660 54350
rect 72156 52780 72212 52836
rect 73276 52220 73332 52276
rect 72044 51548 72100 51604
rect 73276 51602 73332 51604
rect 73276 51550 73278 51602
rect 73278 51550 73330 51602
rect 73330 51550 73332 51602
rect 73276 51548 73332 51550
rect 69804 49810 69860 49812
rect 69804 49758 69806 49810
rect 69806 49758 69858 49810
rect 69858 49758 69860 49810
rect 69804 49756 69860 49758
rect 69244 48636 69300 48692
rect 70140 48242 70196 48244
rect 70140 48190 70142 48242
rect 70142 48190 70194 48242
rect 70194 48190 70196 48242
rect 70140 48188 70196 48190
rect 69244 47346 69300 47348
rect 69244 47294 69246 47346
rect 69246 47294 69298 47346
rect 69298 47294 69300 47346
rect 69244 47292 69300 47294
rect 69020 46620 69076 46676
rect 69692 48130 69748 48132
rect 69692 48078 69694 48130
rect 69694 48078 69746 48130
rect 69746 48078 69748 48130
rect 69692 48076 69748 48078
rect 69804 47234 69860 47236
rect 69804 47182 69806 47234
rect 69806 47182 69858 47234
rect 69858 47182 69860 47234
rect 69804 47180 69860 47182
rect 69356 46396 69412 46452
rect 68796 45052 68852 45108
rect 67900 44268 67956 44324
rect 68460 44098 68516 44100
rect 68460 44046 68462 44098
rect 68462 44046 68514 44098
rect 68514 44046 68516 44098
rect 68460 44044 68516 44046
rect 68236 43762 68292 43764
rect 68236 43710 68238 43762
rect 68238 43710 68290 43762
rect 68290 43710 68292 43762
rect 68236 43708 68292 43710
rect 68460 37772 68516 37828
rect 67564 30044 67620 30100
rect 69356 29932 69412 29988
rect 68124 28588 68180 28644
rect 70364 49644 70420 49700
rect 70364 46620 70420 46676
rect 70812 50092 70868 50148
rect 71708 50316 71764 50372
rect 71932 50092 71988 50148
rect 72156 51378 72212 51380
rect 72156 51326 72158 51378
rect 72158 51326 72210 51378
rect 72210 51326 72212 51378
rect 72156 51324 72212 51326
rect 72380 51378 72436 51380
rect 72380 51326 72382 51378
rect 72382 51326 72434 51378
rect 72434 51326 72436 51378
rect 72380 51324 72436 51326
rect 73500 51324 73556 51380
rect 73724 51100 73780 51156
rect 72268 50428 72324 50484
rect 71484 49756 71540 49812
rect 71148 48748 71204 48804
rect 72268 49922 72324 49924
rect 72268 49870 72270 49922
rect 72270 49870 72322 49922
rect 72322 49870 72324 49922
rect 72268 49868 72324 49870
rect 72268 49698 72324 49700
rect 72268 49646 72270 49698
rect 72270 49646 72322 49698
rect 72322 49646 72324 49698
rect 72268 49644 72324 49646
rect 71484 48748 71540 48804
rect 71372 45500 71428 45556
rect 70252 28588 70308 28644
rect 69356 26460 69412 26516
rect 70812 26012 70868 26068
rect 69468 25788 69524 25844
rect 68796 22092 68852 22148
rect 68796 20524 68852 20580
rect 67788 4450 67844 4452
rect 67788 4398 67790 4450
rect 67790 4398 67842 4450
rect 67842 4398 67844 4450
rect 67788 4396 67844 4398
rect 66780 3724 66836 3780
rect 64092 3388 64148 3444
rect 70588 4396 70644 4452
rect 69132 3388 69188 3444
rect 70476 3442 70532 3444
rect 70476 3390 70478 3442
rect 70478 3390 70530 3442
rect 70530 3390 70532 3442
rect 70476 3388 70532 3390
rect 72268 30098 72324 30100
rect 72268 30046 72270 30098
rect 72270 30046 72322 30098
rect 72322 30046 72324 30098
rect 72268 30044 72324 30046
rect 71372 27692 71428 27748
rect 72716 50316 72772 50372
rect 72492 49868 72548 49924
rect 73164 49868 73220 49924
rect 72380 26012 72436 26068
rect 70924 25788 70980 25844
rect 71820 4450 71876 4452
rect 71820 4398 71822 4450
rect 71822 4398 71874 4450
rect 71874 4398 71876 4450
rect 71820 4396 71876 4398
rect 73724 48748 73780 48804
rect 73276 47570 73332 47572
rect 73276 47518 73278 47570
rect 73278 47518 73330 47570
rect 73330 47518 73332 47570
rect 73276 47516 73332 47518
rect 73276 46844 73332 46900
rect 74172 62466 74228 62468
rect 74172 62414 74174 62466
rect 74174 62414 74226 62466
rect 74226 62414 74228 62466
rect 74172 62412 74228 62414
rect 75628 66274 75684 66276
rect 75628 66222 75630 66274
rect 75630 66222 75682 66274
rect 75682 66222 75684 66274
rect 75628 66220 75684 66222
rect 75180 65324 75236 65380
rect 75852 63420 75908 63476
rect 74508 62300 74564 62356
rect 74732 62354 74788 62356
rect 74732 62302 74734 62354
rect 74734 62302 74786 62354
rect 74786 62302 74788 62354
rect 74732 62300 74788 62302
rect 74508 61682 74564 61684
rect 74508 61630 74510 61682
rect 74510 61630 74562 61682
rect 74562 61630 74564 61682
rect 74508 61628 74564 61630
rect 74172 61180 74228 61236
rect 74060 52274 74116 52276
rect 74060 52222 74062 52274
rect 74062 52222 74114 52274
rect 74114 52222 74116 52274
rect 74060 52220 74116 52222
rect 73948 43372 74004 43428
rect 73948 42812 74004 42868
rect 74060 39564 74116 39620
rect 72716 4172 72772 4228
rect 74060 4226 74116 4228
rect 74060 4174 74062 4226
rect 74062 4174 74114 4226
rect 74114 4174 74116 4226
rect 74060 4172 74116 4174
rect 74956 61346 75012 61348
rect 74956 61294 74958 61346
rect 74958 61294 75010 61346
rect 75010 61294 75012 61346
rect 74956 61292 75012 61294
rect 74284 61010 74340 61012
rect 74284 60958 74286 61010
rect 74286 60958 74338 61010
rect 74338 60958 74340 61010
rect 74284 60956 74340 60958
rect 78988 116562 79044 116564
rect 78988 116510 78990 116562
rect 78990 116510 79042 116562
rect 79042 116510 79044 116562
rect 78988 116508 79044 116510
rect 79772 116508 79828 116564
rect 78764 115724 78820 115780
rect 78988 115778 79044 115780
rect 78988 115726 78990 115778
rect 78990 115726 79042 115778
rect 79042 115726 79044 115778
rect 78988 115724 79044 115726
rect 76524 84866 76580 84868
rect 76524 84814 76526 84866
rect 76526 84814 76578 84866
rect 76578 84814 76580 84866
rect 76524 84812 76580 84814
rect 77084 68796 77140 68852
rect 77868 68796 77924 68852
rect 77644 66892 77700 66948
rect 78316 66892 78372 66948
rect 78876 66332 78932 66388
rect 77420 66220 77476 66276
rect 77196 66162 77252 66164
rect 77196 66110 77198 66162
rect 77198 66110 77250 66162
rect 77250 66110 77252 66162
rect 77196 66108 77252 66110
rect 78204 66108 78260 66164
rect 78428 66220 78484 66276
rect 78428 65548 78484 65604
rect 78652 66220 78708 66276
rect 76412 59948 76468 60004
rect 76636 59948 76692 60004
rect 79548 66386 79604 66388
rect 79548 66334 79550 66386
rect 79550 66334 79602 66386
rect 79602 66334 79604 66386
rect 79548 66332 79604 66334
rect 78652 56364 78708 56420
rect 81564 116562 81620 116564
rect 81564 116510 81566 116562
rect 81566 116510 81618 116562
rect 81618 116510 81620 116562
rect 81564 116508 81620 116510
rect 81228 116284 81284 116340
rect 81276 116058 81332 116060
rect 81276 116006 81278 116058
rect 81278 116006 81330 116058
rect 81330 116006 81332 116058
rect 81276 116004 81332 116006
rect 81380 116058 81436 116060
rect 81380 116006 81382 116058
rect 81382 116006 81434 116058
rect 81434 116006 81436 116058
rect 81380 116004 81436 116006
rect 81484 116058 81540 116060
rect 81484 116006 81486 116058
rect 81486 116006 81538 116058
rect 81538 116006 81540 116058
rect 81484 116004 81540 116006
rect 84812 116956 84868 117012
rect 83468 116508 83524 116564
rect 84812 116562 84868 116564
rect 84812 116510 84814 116562
rect 84814 116510 84866 116562
rect 84866 116510 84868 116562
rect 84812 116508 84868 116510
rect 82572 116338 82628 116340
rect 82572 116286 82574 116338
rect 82574 116286 82626 116338
rect 82626 116286 82628 116338
rect 82572 116284 82628 116286
rect 81900 115724 81956 115780
rect 83244 115778 83300 115780
rect 83244 115726 83246 115778
rect 83246 115726 83298 115778
rect 83298 115726 83300 115778
rect 83244 115724 83300 115726
rect 80444 66892 80500 66948
rect 81276 114490 81332 114492
rect 81276 114438 81278 114490
rect 81278 114438 81330 114490
rect 81330 114438 81332 114490
rect 81276 114436 81332 114438
rect 81380 114490 81436 114492
rect 81380 114438 81382 114490
rect 81382 114438 81434 114490
rect 81434 114438 81436 114490
rect 81380 114436 81436 114438
rect 81484 114490 81540 114492
rect 81484 114438 81486 114490
rect 81486 114438 81538 114490
rect 81538 114438 81540 114490
rect 81484 114436 81540 114438
rect 81276 112922 81332 112924
rect 81276 112870 81278 112922
rect 81278 112870 81330 112922
rect 81330 112870 81332 112922
rect 81276 112868 81332 112870
rect 81380 112922 81436 112924
rect 81380 112870 81382 112922
rect 81382 112870 81434 112922
rect 81434 112870 81436 112922
rect 81380 112868 81436 112870
rect 81484 112922 81540 112924
rect 81484 112870 81486 112922
rect 81486 112870 81538 112922
rect 81538 112870 81540 112922
rect 81484 112868 81540 112870
rect 81276 111354 81332 111356
rect 81276 111302 81278 111354
rect 81278 111302 81330 111354
rect 81330 111302 81332 111354
rect 81276 111300 81332 111302
rect 81380 111354 81436 111356
rect 81380 111302 81382 111354
rect 81382 111302 81434 111354
rect 81434 111302 81436 111354
rect 81380 111300 81436 111302
rect 81484 111354 81540 111356
rect 81484 111302 81486 111354
rect 81486 111302 81538 111354
rect 81538 111302 81540 111354
rect 81484 111300 81540 111302
rect 81276 109786 81332 109788
rect 81276 109734 81278 109786
rect 81278 109734 81330 109786
rect 81330 109734 81332 109786
rect 81276 109732 81332 109734
rect 81380 109786 81436 109788
rect 81380 109734 81382 109786
rect 81382 109734 81434 109786
rect 81434 109734 81436 109786
rect 81380 109732 81436 109734
rect 81484 109786 81540 109788
rect 81484 109734 81486 109786
rect 81486 109734 81538 109786
rect 81538 109734 81540 109786
rect 81484 109732 81540 109734
rect 81276 108218 81332 108220
rect 81276 108166 81278 108218
rect 81278 108166 81330 108218
rect 81330 108166 81332 108218
rect 81276 108164 81332 108166
rect 81380 108218 81436 108220
rect 81380 108166 81382 108218
rect 81382 108166 81434 108218
rect 81434 108166 81436 108218
rect 81380 108164 81436 108166
rect 81484 108218 81540 108220
rect 81484 108166 81486 108218
rect 81486 108166 81538 108218
rect 81538 108166 81540 108218
rect 81484 108164 81540 108166
rect 81276 106650 81332 106652
rect 81276 106598 81278 106650
rect 81278 106598 81330 106650
rect 81330 106598 81332 106650
rect 81276 106596 81332 106598
rect 81380 106650 81436 106652
rect 81380 106598 81382 106650
rect 81382 106598 81434 106650
rect 81434 106598 81436 106650
rect 81380 106596 81436 106598
rect 81484 106650 81540 106652
rect 81484 106598 81486 106650
rect 81486 106598 81538 106650
rect 81538 106598 81540 106650
rect 81484 106596 81540 106598
rect 81276 105082 81332 105084
rect 81276 105030 81278 105082
rect 81278 105030 81330 105082
rect 81330 105030 81332 105082
rect 81276 105028 81332 105030
rect 81380 105082 81436 105084
rect 81380 105030 81382 105082
rect 81382 105030 81434 105082
rect 81434 105030 81436 105082
rect 81380 105028 81436 105030
rect 81484 105082 81540 105084
rect 81484 105030 81486 105082
rect 81486 105030 81538 105082
rect 81538 105030 81540 105082
rect 81484 105028 81540 105030
rect 81276 103514 81332 103516
rect 81276 103462 81278 103514
rect 81278 103462 81330 103514
rect 81330 103462 81332 103514
rect 81276 103460 81332 103462
rect 81380 103514 81436 103516
rect 81380 103462 81382 103514
rect 81382 103462 81434 103514
rect 81434 103462 81436 103514
rect 81380 103460 81436 103462
rect 81484 103514 81540 103516
rect 81484 103462 81486 103514
rect 81486 103462 81538 103514
rect 81538 103462 81540 103514
rect 81484 103460 81540 103462
rect 81276 101946 81332 101948
rect 81276 101894 81278 101946
rect 81278 101894 81330 101946
rect 81330 101894 81332 101946
rect 81276 101892 81332 101894
rect 81380 101946 81436 101948
rect 81380 101894 81382 101946
rect 81382 101894 81434 101946
rect 81434 101894 81436 101946
rect 81380 101892 81436 101894
rect 81484 101946 81540 101948
rect 81484 101894 81486 101946
rect 81486 101894 81538 101946
rect 81538 101894 81540 101946
rect 81484 101892 81540 101894
rect 81276 100378 81332 100380
rect 81276 100326 81278 100378
rect 81278 100326 81330 100378
rect 81330 100326 81332 100378
rect 81276 100324 81332 100326
rect 81380 100378 81436 100380
rect 81380 100326 81382 100378
rect 81382 100326 81434 100378
rect 81434 100326 81436 100378
rect 81380 100324 81436 100326
rect 81484 100378 81540 100380
rect 81484 100326 81486 100378
rect 81486 100326 81538 100378
rect 81538 100326 81540 100378
rect 81484 100324 81540 100326
rect 81276 98810 81332 98812
rect 81276 98758 81278 98810
rect 81278 98758 81330 98810
rect 81330 98758 81332 98810
rect 81276 98756 81332 98758
rect 81380 98810 81436 98812
rect 81380 98758 81382 98810
rect 81382 98758 81434 98810
rect 81434 98758 81436 98810
rect 81380 98756 81436 98758
rect 81484 98810 81540 98812
rect 81484 98758 81486 98810
rect 81486 98758 81538 98810
rect 81538 98758 81540 98810
rect 81484 98756 81540 98758
rect 81276 97242 81332 97244
rect 81276 97190 81278 97242
rect 81278 97190 81330 97242
rect 81330 97190 81332 97242
rect 81276 97188 81332 97190
rect 81380 97242 81436 97244
rect 81380 97190 81382 97242
rect 81382 97190 81434 97242
rect 81434 97190 81436 97242
rect 81380 97188 81436 97190
rect 81484 97242 81540 97244
rect 81484 97190 81486 97242
rect 81486 97190 81538 97242
rect 81538 97190 81540 97242
rect 81484 97188 81540 97190
rect 81276 95674 81332 95676
rect 81276 95622 81278 95674
rect 81278 95622 81330 95674
rect 81330 95622 81332 95674
rect 81276 95620 81332 95622
rect 81380 95674 81436 95676
rect 81380 95622 81382 95674
rect 81382 95622 81434 95674
rect 81434 95622 81436 95674
rect 81380 95620 81436 95622
rect 81484 95674 81540 95676
rect 81484 95622 81486 95674
rect 81486 95622 81538 95674
rect 81538 95622 81540 95674
rect 81484 95620 81540 95622
rect 81276 94106 81332 94108
rect 81276 94054 81278 94106
rect 81278 94054 81330 94106
rect 81330 94054 81332 94106
rect 81276 94052 81332 94054
rect 81380 94106 81436 94108
rect 81380 94054 81382 94106
rect 81382 94054 81434 94106
rect 81434 94054 81436 94106
rect 81380 94052 81436 94054
rect 81484 94106 81540 94108
rect 81484 94054 81486 94106
rect 81486 94054 81538 94106
rect 81538 94054 81540 94106
rect 81484 94052 81540 94054
rect 81276 92538 81332 92540
rect 81276 92486 81278 92538
rect 81278 92486 81330 92538
rect 81330 92486 81332 92538
rect 81276 92484 81332 92486
rect 81380 92538 81436 92540
rect 81380 92486 81382 92538
rect 81382 92486 81434 92538
rect 81434 92486 81436 92538
rect 81380 92484 81436 92486
rect 81484 92538 81540 92540
rect 81484 92486 81486 92538
rect 81486 92486 81538 92538
rect 81538 92486 81540 92538
rect 81484 92484 81540 92486
rect 81276 90970 81332 90972
rect 81276 90918 81278 90970
rect 81278 90918 81330 90970
rect 81330 90918 81332 90970
rect 81276 90916 81332 90918
rect 81380 90970 81436 90972
rect 81380 90918 81382 90970
rect 81382 90918 81434 90970
rect 81434 90918 81436 90970
rect 81380 90916 81436 90918
rect 81484 90970 81540 90972
rect 81484 90918 81486 90970
rect 81486 90918 81538 90970
rect 81538 90918 81540 90970
rect 81484 90916 81540 90918
rect 81276 89402 81332 89404
rect 81276 89350 81278 89402
rect 81278 89350 81330 89402
rect 81330 89350 81332 89402
rect 81276 89348 81332 89350
rect 81380 89402 81436 89404
rect 81380 89350 81382 89402
rect 81382 89350 81434 89402
rect 81434 89350 81436 89402
rect 81380 89348 81436 89350
rect 81484 89402 81540 89404
rect 81484 89350 81486 89402
rect 81486 89350 81538 89402
rect 81538 89350 81540 89402
rect 81484 89348 81540 89350
rect 81276 87834 81332 87836
rect 81276 87782 81278 87834
rect 81278 87782 81330 87834
rect 81330 87782 81332 87834
rect 81276 87780 81332 87782
rect 81380 87834 81436 87836
rect 81380 87782 81382 87834
rect 81382 87782 81434 87834
rect 81434 87782 81436 87834
rect 81380 87780 81436 87782
rect 81484 87834 81540 87836
rect 81484 87782 81486 87834
rect 81486 87782 81538 87834
rect 81538 87782 81540 87834
rect 81484 87780 81540 87782
rect 81276 86266 81332 86268
rect 81276 86214 81278 86266
rect 81278 86214 81330 86266
rect 81330 86214 81332 86266
rect 81276 86212 81332 86214
rect 81380 86266 81436 86268
rect 81380 86214 81382 86266
rect 81382 86214 81434 86266
rect 81434 86214 81436 86266
rect 81380 86212 81436 86214
rect 81484 86266 81540 86268
rect 81484 86214 81486 86266
rect 81486 86214 81538 86266
rect 81538 86214 81540 86266
rect 81484 86212 81540 86214
rect 81276 84698 81332 84700
rect 81276 84646 81278 84698
rect 81278 84646 81330 84698
rect 81330 84646 81332 84698
rect 81276 84644 81332 84646
rect 81380 84698 81436 84700
rect 81380 84646 81382 84698
rect 81382 84646 81434 84698
rect 81434 84646 81436 84698
rect 81380 84644 81436 84646
rect 81484 84698 81540 84700
rect 81484 84646 81486 84698
rect 81486 84646 81538 84698
rect 81538 84646 81540 84698
rect 81484 84644 81540 84646
rect 81276 83130 81332 83132
rect 81276 83078 81278 83130
rect 81278 83078 81330 83130
rect 81330 83078 81332 83130
rect 81276 83076 81332 83078
rect 81380 83130 81436 83132
rect 81380 83078 81382 83130
rect 81382 83078 81434 83130
rect 81434 83078 81436 83130
rect 81380 83076 81436 83078
rect 81484 83130 81540 83132
rect 81484 83078 81486 83130
rect 81486 83078 81538 83130
rect 81538 83078 81540 83130
rect 81484 83076 81540 83078
rect 81276 81562 81332 81564
rect 81276 81510 81278 81562
rect 81278 81510 81330 81562
rect 81330 81510 81332 81562
rect 81276 81508 81332 81510
rect 81380 81562 81436 81564
rect 81380 81510 81382 81562
rect 81382 81510 81434 81562
rect 81434 81510 81436 81562
rect 81380 81508 81436 81510
rect 81484 81562 81540 81564
rect 81484 81510 81486 81562
rect 81486 81510 81538 81562
rect 81538 81510 81540 81562
rect 81484 81508 81540 81510
rect 81276 79994 81332 79996
rect 81276 79942 81278 79994
rect 81278 79942 81330 79994
rect 81330 79942 81332 79994
rect 81276 79940 81332 79942
rect 81380 79994 81436 79996
rect 81380 79942 81382 79994
rect 81382 79942 81434 79994
rect 81434 79942 81436 79994
rect 81380 79940 81436 79942
rect 81484 79994 81540 79996
rect 81484 79942 81486 79994
rect 81486 79942 81538 79994
rect 81538 79942 81540 79994
rect 81484 79940 81540 79942
rect 81276 78426 81332 78428
rect 81276 78374 81278 78426
rect 81278 78374 81330 78426
rect 81330 78374 81332 78426
rect 81276 78372 81332 78374
rect 81380 78426 81436 78428
rect 81380 78374 81382 78426
rect 81382 78374 81434 78426
rect 81434 78374 81436 78426
rect 81380 78372 81436 78374
rect 81484 78426 81540 78428
rect 81484 78374 81486 78426
rect 81486 78374 81538 78426
rect 81538 78374 81540 78426
rect 81484 78372 81540 78374
rect 81276 76858 81332 76860
rect 81276 76806 81278 76858
rect 81278 76806 81330 76858
rect 81330 76806 81332 76858
rect 81276 76804 81332 76806
rect 81380 76858 81436 76860
rect 81380 76806 81382 76858
rect 81382 76806 81434 76858
rect 81434 76806 81436 76858
rect 81380 76804 81436 76806
rect 81484 76858 81540 76860
rect 81484 76806 81486 76858
rect 81486 76806 81538 76858
rect 81538 76806 81540 76858
rect 81484 76804 81540 76806
rect 81276 75290 81332 75292
rect 81276 75238 81278 75290
rect 81278 75238 81330 75290
rect 81330 75238 81332 75290
rect 81276 75236 81332 75238
rect 81380 75290 81436 75292
rect 81380 75238 81382 75290
rect 81382 75238 81434 75290
rect 81434 75238 81436 75290
rect 81380 75236 81436 75238
rect 81484 75290 81540 75292
rect 81484 75238 81486 75290
rect 81486 75238 81538 75290
rect 81538 75238 81540 75290
rect 81484 75236 81540 75238
rect 81276 73722 81332 73724
rect 81276 73670 81278 73722
rect 81278 73670 81330 73722
rect 81330 73670 81332 73722
rect 81276 73668 81332 73670
rect 81380 73722 81436 73724
rect 81380 73670 81382 73722
rect 81382 73670 81434 73722
rect 81434 73670 81436 73722
rect 81380 73668 81436 73670
rect 81484 73722 81540 73724
rect 81484 73670 81486 73722
rect 81486 73670 81538 73722
rect 81538 73670 81540 73722
rect 81484 73668 81540 73670
rect 81276 72154 81332 72156
rect 81276 72102 81278 72154
rect 81278 72102 81330 72154
rect 81330 72102 81332 72154
rect 81276 72100 81332 72102
rect 81380 72154 81436 72156
rect 81380 72102 81382 72154
rect 81382 72102 81434 72154
rect 81434 72102 81436 72154
rect 81380 72100 81436 72102
rect 81484 72154 81540 72156
rect 81484 72102 81486 72154
rect 81486 72102 81538 72154
rect 81538 72102 81540 72154
rect 81484 72100 81540 72102
rect 81276 70586 81332 70588
rect 81276 70534 81278 70586
rect 81278 70534 81330 70586
rect 81330 70534 81332 70586
rect 81276 70532 81332 70534
rect 81380 70586 81436 70588
rect 81380 70534 81382 70586
rect 81382 70534 81434 70586
rect 81434 70534 81436 70586
rect 81380 70532 81436 70534
rect 81484 70586 81540 70588
rect 81484 70534 81486 70586
rect 81486 70534 81538 70586
rect 81538 70534 81540 70586
rect 81484 70532 81540 70534
rect 81276 69018 81332 69020
rect 81276 68966 81278 69018
rect 81278 68966 81330 69018
rect 81330 68966 81332 69018
rect 81276 68964 81332 68966
rect 81380 69018 81436 69020
rect 81380 68966 81382 69018
rect 81382 68966 81434 69018
rect 81434 68966 81436 69018
rect 81380 68964 81436 68966
rect 81484 69018 81540 69020
rect 81484 68966 81486 69018
rect 81486 68966 81538 69018
rect 81538 68966 81540 69018
rect 81484 68964 81540 68966
rect 81276 67450 81332 67452
rect 81276 67398 81278 67450
rect 81278 67398 81330 67450
rect 81330 67398 81332 67450
rect 81276 67396 81332 67398
rect 81380 67450 81436 67452
rect 81380 67398 81382 67450
rect 81382 67398 81434 67450
rect 81434 67398 81436 67450
rect 81380 67396 81436 67398
rect 81484 67450 81540 67452
rect 81484 67398 81486 67450
rect 81486 67398 81538 67450
rect 81538 67398 81540 67450
rect 81484 67396 81540 67398
rect 81228 66946 81284 66948
rect 81228 66894 81230 66946
rect 81230 66894 81282 66946
rect 81282 66894 81284 66946
rect 81228 66892 81284 66894
rect 80556 66332 80612 66388
rect 81676 66050 81732 66052
rect 81676 65998 81678 66050
rect 81678 65998 81730 66050
rect 81730 65998 81732 66050
rect 81676 65996 81732 65998
rect 83132 99820 83188 99876
rect 83132 68012 83188 68068
rect 83244 79324 83300 79380
rect 82348 67282 82404 67284
rect 82348 67230 82350 67282
rect 82350 67230 82402 67282
rect 82402 67230 82404 67282
rect 82348 67228 82404 67230
rect 82236 66220 82292 66276
rect 82012 65996 82068 66052
rect 81276 65882 81332 65884
rect 81276 65830 81278 65882
rect 81278 65830 81330 65882
rect 81330 65830 81332 65882
rect 81276 65828 81332 65830
rect 81380 65882 81436 65884
rect 81380 65830 81382 65882
rect 81382 65830 81434 65882
rect 81434 65830 81436 65882
rect 81380 65828 81436 65830
rect 81484 65882 81540 65884
rect 81484 65830 81486 65882
rect 81486 65830 81538 65882
rect 81538 65830 81540 65882
rect 81484 65828 81540 65830
rect 81276 64314 81332 64316
rect 81276 64262 81278 64314
rect 81278 64262 81330 64314
rect 81330 64262 81332 64314
rect 81276 64260 81332 64262
rect 81380 64314 81436 64316
rect 81380 64262 81382 64314
rect 81382 64262 81434 64314
rect 81434 64262 81436 64314
rect 81380 64260 81436 64262
rect 81484 64314 81540 64316
rect 81484 64262 81486 64314
rect 81486 64262 81538 64314
rect 81538 64262 81540 64314
rect 81484 64260 81540 64262
rect 81276 62746 81332 62748
rect 81276 62694 81278 62746
rect 81278 62694 81330 62746
rect 81330 62694 81332 62746
rect 81276 62692 81332 62694
rect 81380 62746 81436 62748
rect 81380 62694 81382 62746
rect 81382 62694 81434 62746
rect 81434 62694 81436 62746
rect 81380 62692 81436 62694
rect 81484 62746 81540 62748
rect 81484 62694 81486 62746
rect 81486 62694 81538 62746
rect 81538 62694 81540 62746
rect 81484 62692 81540 62694
rect 81116 61570 81172 61572
rect 81116 61518 81118 61570
rect 81118 61518 81170 61570
rect 81170 61518 81172 61570
rect 81116 61516 81172 61518
rect 83020 61570 83076 61572
rect 83020 61518 83022 61570
rect 83022 61518 83074 61570
rect 83074 61518 83076 61570
rect 83020 61516 83076 61518
rect 83356 68012 83412 68068
rect 83356 66444 83412 66500
rect 85260 116396 85316 116452
rect 85932 116450 85988 116452
rect 85932 116398 85934 116450
rect 85934 116398 85986 116450
rect 85986 116398 85988 116450
rect 85932 116396 85988 116398
rect 86604 116956 86660 117012
rect 86156 115836 86212 115892
rect 85260 113372 85316 113428
rect 88172 116508 88228 116564
rect 89068 116562 89124 116564
rect 89068 116510 89070 116562
rect 89070 116510 89122 116562
rect 89122 116510 89124 116562
rect 89068 116508 89124 116510
rect 90860 116508 90916 116564
rect 92652 116562 92708 116564
rect 92652 116510 92654 116562
rect 92654 116510 92706 116562
rect 92706 116510 92708 116562
rect 92652 116508 92708 116510
rect 86940 115836 86996 115892
rect 87948 115666 88004 115668
rect 87948 115614 87950 115666
rect 87950 115614 88002 115666
rect 88002 115614 88004 115666
rect 87948 115612 88004 115614
rect 88284 115612 88340 115668
rect 89852 116396 89908 116452
rect 88172 94556 88228 94612
rect 86268 68124 86324 68180
rect 86492 75628 86548 75684
rect 84140 61628 84196 61684
rect 83244 61404 83300 61460
rect 81276 61178 81332 61180
rect 81276 61126 81278 61178
rect 81278 61126 81330 61178
rect 81330 61126 81332 61178
rect 81276 61124 81332 61126
rect 81380 61178 81436 61180
rect 81380 61126 81382 61178
rect 81382 61126 81434 61178
rect 81434 61126 81436 61178
rect 81380 61124 81436 61126
rect 81484 61178 81540 61180
rect 81484 61126 81486 61178
rect 81486 61126 81538 61178
rect 81538 61126 81540 61178
rect 81484 61124 81540 61126
rect 81276 59610 81332 59612
rect 81276 59558 81278 59610
rect 81278 59558 81330 59610
rect 81330 59558 81332 59610
rect 81276 59556 81332 59558
rect 81380 59610 81436 59612
rect 81380 59558 81382 59610
rect 81382 59558 81434 59610
rect 81434 59558 81436 59610
rect 81380 59556 81436 59558
rect 81484 59610 81540 59612
rect 81484 59558 81486 59610
rect 81486 59558 81538 59610
rect 81538 59558 81540 59610
rect 81484 59556 81540 59558
rect 86492 58716 86548 58772
rect 81276 58042 81332 58044
rect 81276 57990 81278 58042
rect 81278 57990 81330 58042
rect 81330 57990 81332 58042
rect 81276 57988 81332 57990
rect 81380 58042 81436 58044
rect 81380 57990 81382 58042
rect 81382 57990 81434 58042
rect 81434 57990 81436 58042
rect 81380 57988 81436 57990
rect 81484 58042 81540 58044
rect 81484 57990 81486 58042
rect 81486 57990 81538 58042
rect 81538 57990 81540 58042
rect 81484 57988 81540 57990
rect 83132 57820 83188 57876
rect 79772 56252 79828 56308
rect 80108 56924 80164 56980
rect 76636 54572 76692 54628
rect 79436 54460 79492 54516
rect 77868 53340 77924 53396
rect 76972 50652 77028 50708
rect 76972 48748 77028 48804
rect 75068 43372 75124 43428
rect 75068 29986 75124 29988
rect 75068 29934 75070 29986
rect 75070 29934 75122 29986
rect 75122 29934 75124 29986
rect 75068 29932 75124 29934
rect 76524 30044 76580 30100
rect 76524 22316 76580 22372
rect 79772 44380 79828 44436
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 80332 56194 80388 56196
rect 80332 56142 80334 56194
rect 80334 56142 80386 56194
rect 80386 56142 80388 56194
rect 80332 56140 80388 56142
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 80556 48076 80612 48132
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 80556 44828 80612 44884
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 82348 43426 82404 43428
rect 82348 43374 82350 43426
rect 82350 43374 82402 43426
rect 82402 43374 82404 43426
rect 82348 43372 82404 43374
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 80108 26236 80164 26292
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 79772 24892 79828 24948
rect 78316 23714 78372 23716
rect 78316 23662 78318 23714
rect 78318 23662 78370 23714
rect 78370 23662 78372 23714
rect 78316 23660 78372 23662
rect 77644 23154 77700 23156
rect 77644 23102 77646 23154
rect 77646 23102 77698 23154
rect 77698 23102 77700 23154
rect 77644 23100 77700 23102
rect 78540 23154 78596 23156
rect 78540 23102 78542 23154
rect 78542 23102 78594 23154
rect 78594 23102 78596 23154
rect 78540 23100 78596 23102
rect 79100 23660 79156 23716
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 77532 22370 77588 22372
rect 77532 22318 77534 22370
rect 77534 22318 77586 22370
rect 77586 22318 77588 22370
rect 77532 22316 77588 22318
rect 77532 21420 77588 21476
rect 74060 3388 74116 3444
rect 75068 3442 75124 3444
rect 75068 3390 75070 3442
rect 75070 3390 75122 3442
rect 75122 3390 75124 3442
rect 75068 3388 75124 3390
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 88172 55692 88228 55748
rect 88508 58380 88564 58436
rect 96636 116842 96692 116844
rect 96636 116790 96638 116842
rect 96638 116790 96690 116842
rect 96690 116790 96692 116842
rect 96636 116788 96692 116790
rect 96740 116842 96796 116844
rect 96740 116790 96742 116842
rect 96742 116790 96794 116842
rect 96794 116790 96796 116842
rect 96740 116788 96796 116790
rect 96844 116842 96900 116844
rect 96844 116790 96846 116842
rect 96846 116790 96898 116842
rect 96898 116790 96900 116842
rect 96844 116788 96900 116790
rect 95900 116396 95956 116452
rect 95116 116284 95172 116340
rect 96908 116338 96964 116340
rect 96908 116286 96910 116338
rect 96910 116286 96962 116338
rect 96962 116286 96964 116338
rect 96908 116284 96964 116286
rect 99372 116284 99428 116340
rect 96636 115274 96692 115276
rect 96636 115222 96638 115274
rect 96638 115222 96690 115274
rect 96690 115222 96692 115274
rect 96636 115220 96692 115222
rect 96740 115274 96796 115276
rect 96740 115222 96742 115274
rect 96742 115222 96794 115274
rect 96794 115222 96796 115274
rect 96740 115220 96796 115222
rect 96844 115274 96900 115276
rect 96844 115222 96846 115274
rect 96846 115222 96898 115274
rect 96898 115222 96900 115274
rect 96844 115220 96900 115222
rect 96636 113706 96692 113708
rect 96636 113654 96638 113706
rect 96638 113654 96690 113706
rect 96690 113654 96692 113706
rect 96636 113652 96692 113654
rect 96740 113706 96796 113708
rect 96740 113654 96742 113706
rect 96742 113654 96794 113706
rect 96794 113654 96796 113706
rect 96740 113652 96796 113654
rect 96844 113706 96900 113708
rect 96844 113654 96846 113706
rect 96846 113654 96898 113706
rect 96898 113654 96900 113706
rect 96844 113652 96900 113654
rect 96636 112138 96692 112140
rect 96636 112086 96638 112138
rect 96638 112086 96690 112138
rect 96690 112086 96692 112138
rect 96636 112084 96692 112086
rect 96740 112138 96796 112140
rect 96740 112086 96742 112138
rect 96742 112086 96794 112138
rect 96794 112086 96796 112138
rect 96740 112084 96796 112086
rect 96844 112138 96900 112140
rect 96844 112086 96846 112138
rect 96846 112086 96898 112138
rect 96898 112086 96900 112138
rect 96844 112084 96900 112086
rect 96636 110570 96692 110572
rect 96636 110518 96638 110570
rect 96638 110518 96690 110570
rect 96690 110518 96692 110570
rect 96636 110516 96692 110518
rect 96740 110570 96796 110572
rect 96740 110518 96742 110570
rect 96742 110518 96794 110570
rect 96794 110518 96796 110570
rect 96740 110516 96796 110518
rect 96844 110570 96900 110572
rect 96844 110518 96846 110570
rect 96846 110518 96898 110570
rect 96898 110518 96900 110570
rect 96844 110516 96900 110518
rect 91196 68012 91252 68068
rect 93212 109228 93268 109284
rect 89852 57484 89908 57540
rect 91532 64652 91588 64708
rect 89964 54626 90020 54628
rect 89964 54574 89966 54626
rect 89966 54574 90018 54626
rect 90018 54574 90020 54626
rect 89964 54572 90020 54574
rect 88508 54460 88564 54516
rect 84812 54348 84868 54404
rect 83132 5852 83188 5908
rect 84140 27692 84196 27748
rect 81676 4844 81732 4900
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 78316 4284 78372 4340
rect 78876 4338 78932 4340
rect 78876 4286 78878 4338
rect 78878 4286 78930 4338
rect 78930 4286 78932 4338
rect 78876 4284 78932 4286
rect 78764 4172 78820 4228
rect 75740 3388 75796 3444
rect 75404 3276 75460 3332
rect 76300 3330 76356 3332
rect 76300 3278 76302 3330
rect 76302 3278 76354 3330
rect 76354 3278 76356 3330
rect 76300 3276 76356 3278
rect 79548 4226 79604 4228
rect 79548 4174 79550 4226
rect 79550 4174 79602 4226
rect 79602 4174 79604 4226
rect 79548 4172 79604 4174
rect 81676 4562 81732 4564
rect 81676 4510 81678 4562
rect 81678 4510 81730 4562
rect 81730 4510 81732 4562
rect 81676 4508 81732 4510
rect 83468 4508 83524 4564
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 89628 54514 89684 54516
rect 89628 54462 89630 54514
rect 89630 54462 89682 54514
rect 89682 54462 89684 54514
rect 89628 54460 89684 54462
rect 86492 47404 86548 47460
rect 87276 43372 87332 43428
rect 87836 43426 87892 43428
rect 87836 43374 87838 43426
rect 87838 43374 87890 43426
rect 87890 43374 87892 43426
rect 87836 43372 87892 43374
rect 86492 24444 86548 24500
rect 86940 24892 86996 24948
rect 84812 17612 84868 17668
rect 86604 4396 86660 4452
rect 83468 3442 83524 3444
rect 83468 3390 83470 3442
rect 83470 3390 83522 3442
rect 83522 3390 83524 3442
rect 83468 3388 83524 3390
rect 85148 3442 85204 3444
rect 85148 3390 85150 3442
rect 85150 3390 85202 3442
rect 85202 3390 85204 3442
rect 85148 3388 85204 3390
rect 87948 4450 88004 4452
rect 87948 4398 87950 4450
rect 87950 4398 88002 4450
rect 88002 4398 88004 4450
rect 87948 4396 88004 4398
rect 96636 109002 96692 109004
rect 96636 108950 96638 109002
rect 96638 108950 96690 109002
rect 96690 108950 96692 109002
rect 96636 108948 96692 108950
rect 96740 109002 96796 109004
rect 96740 108950 96742 109002
rect 96742 108950 96794 109002
rect 96794 108950 96796 109002
rect 96740 108948 96796 108950
rect 96844 109002 96900 109004
rect 96844 108950 96846 109002
rect 96846 108950 96898 109002
rect 96898 108950 96900 109002
rect 96844 108948 96900 108950
rect 96636 107434 96692 107436
rect 96636 107382 96638 107434
rect 96638 107382 96690 107434
rect 96690 107382 96692 107434
rect 96636 107380 96692 107382
rect 96740 107434 96796 107436
rect 96740 107382 96742 107434
rect 96742 107382 96794 107434
rect 96794 107382 96796 107434
rect 96740 107380 96796 107382
rect 96844 107434 96900 107436
rect 96844 107382 96846 107434
rect 96846 107382 96898 107434
rect 96898 107382 96900 107434
rect 96844 107380 96900 107382
rect 96636 105866 96692 105868
rect 96636 105814 96638 105866
rect 96638 105814 96690 105866
rect 96690 105814 96692 105866
rect 96636 105812 96692 105814
rect 96740 105866 96796 105868
rect 96740 105814 96742 105866
rect 96742 105814 96794 105866
rect 96794 105814 96796 105866
rect 96740 105812 96796 105814
rect 96844 105866 96900 105868
rect 96844 105814 96846 105866
rect 96846 105814 96898 105866
rect 96898 105814 96900 105866
rect 96844 105812 96900 105814
rect 100828 116338 100884 116340
rect 100828 116286 100830 116338
rect 100830 116286 100882 116338
rect 100882 116286 100884 116338
rect 100828 116284 100884 116286
rect 101612 116508 101668 116564
rect 100940 115500 100996 115556
rect 100492 115388 100548 115444
rect 101052 115388 101108 115444
rect 99820 105196 99876 105252
rect 100044 104524 100100 104580
rect 96636 104298 96692 104300
rect 96636 104246 96638 104298
rect 96638 104246 96690 104298
rect 96690 104246 96692 104298
rect 96636 104244 96692 104246
rect 96740 104298 96796 104300
rect 96740 104246 96742 104298
rect 96742 104246 96794 104298
rect 96794 104246 96796 104298
rect 96740 104244 96796 104246
rect 96844 104298 96900 104300
rect 96844 104246 96846 104298
rect 96846 104246 96898 104298
rect 96898 104246 96900 104298
rect 96844 104244 96900 104246
rect 96636 102730 96692 102732
rect 96636 102678 96638 102730
rect 96638 102678 96690 102730
rect 96690 102678 96692 102730
rect 96636 102676 96692 102678
rect 96740 102730 96796 102732
rect 96740 102678 96742 102730
rect 96742 102678 96794 102730
rect 96794 102678 96796 102730
rect 96740 102676 96796 102678
rect 96844 102730 96900 102732
rect 96844 102678 96846 102730
rect 96846 102678 96898 102730
rect 96898 102678 96900 102730
rect 96844 102676 96900 102678
rect 96636 101162 96692 101164
rect 96636 101110 96638 101162
rect 96638 101110 96690 101162
rect 96690 101110 96692 101162
rect 96636 101108 96692 101110
rect 96740 101162 96796 101164
rect 96740 101110 96742 101162
rect 96742 101110 96794 101162
rect 96794 101110 96796 101162
rect 96740 101108 96796 101110
rect 96844 101162 96900 101164
rect 96844 101110 96846 101162
rect 96846 101110 96898 101162
rect 96898 101110 96900 101162
rect 96844 101108 96900 101110
rect 96636 99594 96692 99596
rect 96636 99542 96638 99594
rect 96638 99542 96690 99594
rect 96690 99542 96692 99594
rect 96636 99540 96692 99542
rect 96740 99594 96796 99596
rect 96740 99542 96742 99594
rect 96742 99542 96794 99594
rect 96794 99542 96796 99594
rect 96740 99540 96796 99542
rect 96844 99594 96900 99596
rect 96844 99542 96846 99594
rect 96846 99542 96898 99594
rect 96898 99542 96900 99594
rect 96844 99540 96900 99542
rect 96636 98026 96692 98028
rect 96636 97974 96638 98026
rect 96638 97974 96690 98026
rect 96690 97974 96692 98026
rect 96636 97972 96692 97974
rect 96740 98026 96796 98028
rect 96740 97974 96742 98026
rect 96742 97974 96794 98026
rect 96794 97974 96796 98026
rect 96740 97972 96796 97974
rect 96844 98026 96900 98028
rect 96844 97974 96846 98026
rect 96846 97974 96898 98026
rect 96898 97974 96900 98026
rect 96844 97972 96900 97974
rect 96636 96458 96692 96460
rect 96636 96406 96638 96458
rect 96638 96406 96690 96458
rect 96690 96406 96692 96458
rect 96636 96404 96692 96406
rect 96740 96458 96796 96460
rect 96740 96406 96742 96458
rect 96742 96406 96794 96458
rect 96794 96406 96796 96458
rect 96740 96404 96796 96406
rect 96844 96458 96900 96460
rect 96844 96406 96846 96458
rect 96846 96406 96898 96458
rect 96898 96406 96900 96458
rect 96844 96404 96900 96406
rect 96636 94890 96692 94892
rect 96636 94838 96638 94890
rect 96638 94838 96690 94890
rect 96690 94838 96692 94890
rect 96636 94836 96692 94838
rect 96740 94890 96796 94892
rect 96740 94838 96742 94890
rect 96742 94838 96794 94890
rect 96794 94838 96796 94890
rect 96740 94836 96796 94838
rect 96844 94890 96900 94892
rect 96844 94838 96846 94890
rect 96846 94838 96898 94890
rect 96898 94838 96900 94890
rect 96844 94836 96900 94838
rect 96636 93322 96692 93324
rect 96636 93270 96638 93322
rect 96638 93270 96690 93322
rect 96690 93270 96692 93322
rect 96636 93268 96692 93270
rect 96740 93322 96796 93324
rect 96740 93270 96742 93322
rect 96742 93270 96794 93322
rect 96794 93270 96796 93322
rect 96740 93268 96796 93270
rect 96844 93322 96900 93324
rect 96844 93270 96846 93322
rect 96846 93270 96898 93322
rect 96898 93270 96900 93322
rect 96844 93268 96900 93270
rect 98252 92876 98308 92932
rect 96636 91754 96692 91756
rect 96636 91702 96638 91754
rect 96638 91702 96690 91754
rect 96690 91702 96692 91754
rect 96636 91700 96692 91702
rect 96740 91754 96796 91756
rect 96740 91702 96742 91754
rect 96742 91702 96794 91754
rect 96794 91702 96796 91754
rect 96740 91700 96796 91702
rect 96844 91754 96900 91756
rect 96844 91702 96846 91754
rect 96846 91702 96898 91754
rect 96898 91702 96900 91754
rect 96844 91700 96900 91702
rect 96636 90186 96692 90188
rect 96636 90134 96638 90186
rect 96638 90134 96690 90186
rect 96690 90134 96692 90186
rect 96636 90132 96692 90134
rect 96740 90186 96796 90188
rect 96740 90134 96742 90186
rect 96742 90134 96794 90186
rect 96794 90134 96796 90186
rect 96740 90132 96796 90134
rect 96844 90186 96900 90188
rect 96844 90134 96846 90186
rect 96846 90134 96898 90186
rect 96898 90134 96900 90186
rect 96844 90132 96900 90134
rect 96636 88618 96692 88620
rect 96636 88566 96638 88618
rect 96638 88566 96690 88618
rect 96690 88566 96692 88618
rect 96636 88564 96692 88566
rect 96740 88618 96796 88620
rect 96740 88566 96742 88618
rect 96742 88566 96794 88618
rect 96794 88566 96796 88618
rect 96740 88564 96796 88566
rect 96844 88618 96900 88620
rect 96844 88566 96846 88618
rect 96846 88566 96898 88618
rect 96898 88566 96900 88618
rect 96844 88564 96900 88566
rect 96636 87050 96692 87052
rect 96636 86998 96638 87050
rect 96638 86998 96690 87050
rect 96690 86998 96692 87050
rect 96636 86996 96692 86998
rect 96740 87050 96796 87052
rect 96740 86998 96742 87050
rect 96742 86998 96794 87050
rect 96794 86998 96796 87050
rect 96740 86996 96796 86998
rect 96844 87050 96900 87052
rect 96844 86998 96846 87050
rect 96846 86998 96898 87050
rect 96898 86998 96900 87050
rect 96844 86996 96900 86998
rect 96636 85482 96692 85484
rect 96636 85430 96638 85482
rect 96638 85430 96690 85482
rect 96690 85430 96692 85482
rect 96636 85428 96692 85430
rect 96740 85482 96796 85484
rect 96740 85430 96742 85482
rect 96742 85430 96794 85482
rect 96794 85430 96796 85482
rect 96740 85428 96796 85430
rect 96844 85482 96900 85484
rect 96844 85430 96846 85482
rect 96846 85430 96898 85482
rect 96898 85430 96900 85482
rect 96844 85428 96900 85430
rect 96636 83914 96692 83916
rect 96636 83862 96638 83914
rect 96638 83862 96690 83914
rect 96690 83862 96692 83914
rect 96636 83860 96692 83862
rect 96740 83914 96796 83916
rect 96740 83862 96742 83914
rect 96742 83862 96794 83914
rect 96794 83862 96796 83914
rect 96740 83860 96796 83862
rect 96844 83914 96900 83916
rect 96844 83862 96846 83914
rect 96846 83862 96898 83914
rect 96898 83862 96900 83914
rect 96844 83860 96900 83862
rect 96636 82346 96692 82348
rect 96636 82294 96638 82346
rect 96638 82294 96690 82346
rect 96690 82294 96692 82346
rect 96636 82292 96692 82294
rect 96740 82346 96796 82348
rect 96740 82294 96742 82346
rect 96742 82294 96794 82346
rect 96794 82294 96796 82346
rect 96740 82292 96796 82294
rect 96844 82346 96900 82348
rect 96844 82294 96846 82346
rect 96846 82294 96898 82346
rect 96898 82294 96900 82346
rect 96844 82292 96900 82294
rect 96636 80778 96692 80780
rect 96636 80726 96638 80778
rect 96638 80726 96690 80778
rect 96690 80726 96692 80778
rect 96636 80724 96692 80726
rect 96740 80778 96796 80780
rect 96740 80726 96742 80778
rect 96742 80726 96794 80778
rect 96794 80726 96796 80778
rect 96740 80724 96796 80726
rect 96844 80778 96900 80780
rect 96844 80726 96846 80778
rect 96846 80726 96898 80778
rect 96898 80726 96900 80778
rect 96844 80724 96900 80726
rect 96636 79210 96692 79212
rect 96636 79158 96638 79210
rect 96638 79158 96690 79210
rect 96690 79158 96692 79210
rect 96636 79156 96692 79158
rect 96740 79210 96796 79212
rect 96740 79158 96742 79210
rect 96742 79158 96794 79210
rect 96794 79158 96796 79210
rect 96740 79156 96796 79158
rect 96844 79210 96900 79212
rect 96844 79158 96846 79210
rect 96846 79158 96898 79210
rect 96898 79158 96900 79210
rect 96844 79156 96900 79158
rect 96636 77642 96692 77644
rect 96636 77590 96638 77642
rect 96638 77590 96690 77642
rect 96690 77590 96692 77642
rect 96636 77588 96692 77590
rect 96740 77642 96796 77644
rect 96740 77590 96742 77642
rect 96742 77590 96794 77642
rect 96794 77590 96796 77642
rect 96740 77588 96796 77590
rect 96844 77642 96900 77644
rect 96844 77590 96846 77642
rect 96846 77590 96898 77642
rect 96898 77590 96900 77642
rect 96844 77588 96900 77590
rect 96636 76074 96692 76076
rect 96636 76022 96638 76074
rect 96638 76022 96690 76074
rect 96690 76022 96692 76074
rect 96636 76020 96692 76022
rect 96740 76074 96796 76076
rect 96740 76022 96742 76074
rect 96742 76022 96794 76074
rect 96794 76022 96796 76074
rect 96740 76020 96796 76022
rect 96844 76074 96900 76076
rect 96844 76022 96846 76074
rect 96846 76022 96898 76074
rect 96898 76022 96900 76074
rect 96844 76020 96900 76022
rect 96636 74506 96692 74508
rect 96636 74454 96638 74506
rect 96638 74454 96690 74506
rect 96690 74454 96692 74506
rect 96636 74452 96692 74454
rect 96740 74506 96796 74508
rect 96740 74454 96742 74506
rect 96742 74454 96794 74506
rect 96794 74454 96796 74506
rect 96740 74452 96796 74454
rect 96844 74506 96900 74508
rect 96844 74454 96846 74506
rect 96846 74454 96898 74506
rect 96898 74454 96900 74506
rect 96844 74452 96900 74454
rect 96636 72938 96692 72940
rect 96636 72886 96638 72938
rect 96638 72886 96690 72938
rect 96690 72886 96692 72938
rect 96636 72884 96692 72886
rect 96740 72938 96796 72940
rect 96740 72886 96742 72938
rect 96742 72886 96794 72938
rect 96794 72886 96796 72938
rect 96740 72884 96796 72886
rect 96844 72938 96900 72940
rect 96844 72886 96846 72938
rect 96846 72886 96898 72938
rect 96898 72886 96900 72938
rect 96844 72884 96900 72886
rect 96636 71370 96692 71372
rect 96636 71318 96638 71370
rect 96638 71318 96690 71370
rect 96690 71318 96692 71370
rect 96636 71316 96692 71318
rect 96740 71370 96796 71372
rect 96740 71318 96742 71370
rect 96742 71318 96794 71370
rect 96794 71318 96796 71370
rect 96740 71316 96796 71318
rect 96844 71370 96900 71372
rect 96844 71318 96846 71370
rect 96846 71318 96898 71370
rect 96898 71318 96900 71370
rect 96844 71316 96900 71318
rect 96636 69802 96692 69804
rect 96636 69750 96638 69802
rect 96638 69750 96690 69802
rect 96690 69750 96692 69802
rect 96636 69748 96692 69750
rect 96740 69802 96796 69804
rect 96740 69750 96742 69802
rect 96742 69750 96794 69802
rect 96794 69750 96796 69802
rect 96740 69748 96796 69750
rect 96844 69802 96900 69804
rect 96844 69750 96846 69802
rect 96846 69750 96898 69802
rect 96898 69750 96900 69802
rect 96844 69748 96900 69750
rect 96636 68234 96692 68236
rect 96636 68182 96638 68234
rect 96638 68182 96690 68234
rect 96690 68182 96692 68234
rect 96636 68180 96692 68182
rect 96740 68234 96796 68236
rect 96740 68182 96742 68234
rect 96742 68182 96794 68234
rect 96794 68182 96796 68234
rect 96740 68180 96796 68182
rect 96844 68234 96900 68236
rect 96844 68182 96846 68234
rect 96846 68182 96898 68234
rect 96898 68182 96900 68234
rect 96844 68180 96900 68182
rect 96636 66666 96692 66668
rect 96636 66614 96638 66666
rect 96638 66614 96690 66666
rect 96690 66614 96692 66666
rect 96636 66612 96692 66614
rect 96740 66666 96796 66668
rect 96740 66614 96742 66666
rect 96742 66614 96794 66666
rect 96794 66614 96796 66666
rect 96740 66612 96796 66614
rect 96844 66666 96900 66668
rect 96844 66614 96846 66666
rect 96846 66614 96898 66666
rect 96898 66614 96900 66666
rect 96844 66612 96900 66614
rect 96636 65098 96692 65100
rect 96636 65046 96638 65098
rect 96638 65046 96690 65098
rect 96690 65046 96692 65098
rect 96636 65044 96692 65046
rect 96740 65098 96796 65100
rect 96740 65046 96742 65098
rect 96742 65046 96794 65098
rect 96794 65046 96796 65098
rect 96740 65044 96796 65046
rect 96844 65098 96900 65100
rect 96844 65046 96846 65098
rect 96846 65046 96898 65098
rect 96898 65046 96900 65098
rect 96844 65044 96900 65046
rect 96636 63530 96692 63532
rect 96636 63478 96638 63530
rect 96638 63478 96690 63530
rect 96690 63478 96692 63530
rect 96636 63476 96692 63478
rect 96740 63530 96796 63532
rect 96740 63478 96742 63530
rect 96742 63478 96794 63530
rect 96794 63478 96796 63530
rect 96740 63476 96796 63478
rect 96844 63530 96900 63532
rect 96844 63478 96846 63530
rect 96846 63478 96898 63530
rect 96898 63478 96900 63530
rect 96844 63476 96900 63478
rect 98252 62300 98308 62356
rect 96636 61962 96692 61964
rect 96636 61910 96638 61962
rect 96638 61910 96690 61962
rect 96690 61910 96692 61962
rect 96636 61908 96692 61910
rect 96740 61962 96796 61964
rect 96740 61910 96742 61962
rect 96742 61910 96794 61962
rect 96794 61910 96796 61962
rect 96740 61908 96796 61910
rect 96844 61962 96900 61964
rect 96844 61910 96846 61962
rect 96846 61910 96898 61962
rect 96898 61910 96900 61962
rect 96844 61908 96900 61910
rect 98252 61740 98308 61796
rect 96636 60394 96692 60396
rect 96636 60342 96638 60394
rect 96638 60342 96690 60394
rect 96690 60342 96692 60394
rect 96636 60340 96692 60342
rect 96740 60394 96796 60396
rect 96740 60342 96742 60394
rect 96742 60342 96794 60394
rect 96794 60342 96796 60394
rect 96740 60340 96796 60342
rect 96844 60394 96900 60396
rect 96844 60342 96846 60394
rect 96846 60342 96898 60394
rect 96898 60342 96900 60394
rect 96844 60340 96900 60342
rect 96636 58826 96692 58828
rect 96636 58774 96638 58826
rect 96638 58774 96690 58826
rect 96690 58774 96692 58826
rect 96636 58772 96692 58774
rect 96740 58826 96796 58828
rect 96740 58774 96742 58826
rect 96742 58774 96794 58826
rect 96794 58774 96796 58826
rect 96740 58772 96796 58774
rect 96844 58826 96900 58828
rect 96844 58774 96846 58826
rect 96846 58774 96898 58826
rect 96898 58774 96900 58826
rect 96844 58772 96900 58774
rect 96636 57258 96692 57260
rect 96636 57206 96638 57258
rect 96638 57206 96690 57258
rect 96690 57206 96692 57258
rect 96636 57204 96692 57206
rect 96740 57258 96796 57260
rect 96740 57206 96742 57258
rect 96742 57206 96794 57258
rect 96794 57206 96796 57258
rect 96740 57204 96796 57206
rect 96844 57258 96900 57260
rect 96844 57206 96846 57258
rect 96846 57206 96898 57258
rect 96898 57206 96900 57258
rect 96844 57204 96900 57206
rect 93212 55804 93268 55860
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 91532 51324 91588 51380
rect 92988 54684 93044 54740
rect 90188 50428 90244 50484
rect 90076 20578 90132 20580
rect 90076 20526 90078 20578
rect 90078 20526 90130 20578
rect 90130 20526 90132 20578
rect 90076 20524 90132 20526
rect 91532 47516 91588 47572
rect 91532 41916 91588 41972
rect 91868 40908 91924 40964
rect 90636 21474 90692 21476
rect 90636 21422 90638 21474
rect 90638 21422 90690 21474
rect 90690 21422 90692 21474
rect 90636 21420 90692 21422
rect 91308 21586 91364 21588
rect 91308 21534 91310 21586
rect 91310 21534 91362 21586
rect 91362 21534 91364 21586
rect 91308 21532 91364 21534
rect 90524 20748 90580 20804
rect 91532 20802 91588 20804
rect 91532 20750 91534 20802
rect 91534 20750 91586 20802
rect 91586 20750 91588 20802
rect 91532 20748 91588 20750
rect 92204 20802 92260 20804
rect 92204 20750 92206 20802
rect 92206 20750 92258 20802
rect 92258 20750 92260 20802
rect 92204 20748 92260 20750
rect 92316 20690 92372 20692
rect 92316 20638 92318 20690
rect 92318 20638 92370 20690
rect 92370 20638 92372 20690
rect 92316 20636 92372 20638
rect 92204 20524 92260 20580
rect 90524 4508 90580 4564
rect 90188 4284 90244 4340
rect 92652 4396 92708 4452
rect 88508 3500 88564 3556
rect 89964 3554 90020 3556
rect 89964 3502 89966 3554
rect 89966 3502 90018 3554
rect 90018 3502 90020 3554
rect 89964 3500 90020 3502
rect 91308 3442 91364 3444
rect 91308 3390 91310 3442
rect 91310 3390 91362 3442
rect 91362 3390 91364 3442
rect 91308 3388 91364 3390
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 96636 47850 96692 47852
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 96636 46282 96692 46284
rect 94892 46172 94948 46228
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 95676 35644 95732 35700
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 95676 34636 95732 34692
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 94892 33516 94948 33572
rect 95228 32396 95284 32452
rect 93100 21420 93156 21476
rect 94108 21474 94164 21476
rect 94108 21422 94110 21474
rect 94110 21422 94162 21474
rect 94162 21422 94164 21474
rect 94108 21420 94164 21422
rect 95004 21420 95060 21476
rect 93100 20636 93156 20692
rect 93996 4450 94052 4452
rect 93996 4398 93998 4450
rect 93998 4398 94050 4450
rect 94050 4398 94052 4450
rect 93996 4396 94052 4398
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 95228 20748 95284 20804
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 106876 116284 106932 116340
rect 101724 115554 101780 115556
rect 101724 115502 101726 115554
rect 101726 115502 101778 115554
rect 101778 115502 101780 115554
rect 101724 115500 101780 115502
rect 103292 115500 103348 115556
rect 106652 107660 106708 107716
rect 103292 62524 103348 62580
rect 104972 74172 105028 74228
rect 103516 55468 103572 55524
rect 101612 54236 101668 54292
rect 101836 55244 101892 55300
rect 100044 51996 100100 52052
rect 100268 51100 100324 51156
rect 100828 43372 100884 43428
rect 101836 43372 101892 43428
rect 100828 41132 100884 41188
rect 100268 14252 100324 14308
rect 101836 40348 101892 40404
rect 101836 12012 101892 12068
rect 103292 37772 103348 37828
rect 98252 6748 98308 6804
rect 100268 9212 100324 9268
rect 96348 5852 96404 5908
rect 92988 3442 93044 3444
rect 92988 3390 92990 3442
rect 92990 3390 93042 3442
rect 93042 3390 93044 3442
rect 92988 3388 93044 3390
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 99148 5010 99204 5012
rect 99148 4958 99150 5010
rect 99150 4958 99202 5010
rect 99202 4958 99204 5010
rect 99148 4956 99204 4958
rect 99932 4956 99988 5012
rect 98028 4396 98084 4452
rect 99372 4450 99428 4452
rect 99372 4398 99374 4450
rect 99374 4398 99426 4450
rect 99426 4398 99428 4450
rect 99372 4396 99428 4398
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 96012 3388 96068 3444
rect 97356 3442 97412 3444
rect 97356 3390 97358 3442
rect 97358 3390 97410 3442
rect 97410 3390 97412 3442
rect 97356 3388 97412 3390
rect 98364 4284 98420 4340
rect 99932 4284 99988 4340
rect 101388 4508 101444 4564
rect 108668 116338 108724 116340
rect 108668 116286 108670 116338
rect 108670 116286 108722 116338
rect 108722 116286 108724 116338
rect 108668 116284 108724 116286
rect 108780 115724 108836 115780
rect 110124 115778 110180 115780
rect 110124 115726 110126 115778
rect 110126 115726 110178 115778
rect 110178 115726 110180 115778
rect 110124 115724 110180 115726
rect 111804 116562 111860 116564
rect 111804 116510 111806 116562
rect 111806 116510 111858 116562
rect 111858 116510 111860 116562
rect 111804 116508 111860 116510
rect 110908 116284 110964 116340
rect 112812 116338 112868 116340
rect 112812 116286 112814 116338
rect 112814 116286 112866 116338
rect 112866 116286 112868 116338
rect 112812 116284 112868 116286
rect 115724 116562 115780 116564
rect 115724 116510 115726 116562
rect 115726 116510 115778 116562
rect 115778 116510 115780 116562
rect 115724 116508 115780 116510
rect 114828 116284 114884 116340
rect 116508 116338 116564 116340
rect 116508 116286 116510 116338
rect 116510 116286 116562 116338
rect 116562 116286 116564 116338
rect 116508 116284 116564 116286
rect 111996 116058 112052 116060
rect 111996 116006 111998 116058
rect 111998 116006 112050 116058
rect 112050 116006 112052 116058
rect 111996 116004 112052 116006
rect 112100 116058 112156 116060
rect 112100 116006 112102 116058
rect 112102 116006 112154 116058
rect 112154 116006 112156 116058
rect 112100 116004 112156 116006
rect 112204 116058 112260 116060
rect 112204 116006 112206 116058
rect 112206 116006 112258 116058
rect 112258 116006 112260 116058
rect 112204 116004 112260 116006
rect 110348 115724 110404 115780
rect 111244 115778 111300 115780
rect 111244 115726 111246 115778
rect 111246 115726 111298 115778
rect 111298 115726 111300 115778
rect 111244 115724 111300 115726
rect 109116 115554 109172 115556
rect 109116 115502 109118 115554
rect 109118 115502 109170 115554
rect 109170 115502 109172 115554
rect 109116 115500 109172 115502
rect 110796 114882 110852 114884
rect 110796 114830 110798 114882
rect 110798 114830 110850 114882
rect 110850 114830 110852 114882
rect 110796 114828 110852 114830
rect 115500 115554 115556 115556
rect 115500 115502 115502 115554
rect 115502 115502 115554 115554
rect 115554 115502 115556 115554
rect 115500 115500 115556 115502
rect 115836 115276 115892 115332
rect 115500 115164 115556 115220
rect 112588 114828 112644 114884
rect 111996 114490 112052 114492
rect 111996 114438 111998 114490
rect 111998 114438 112050 114490
rect 112050 114438 112052 114490
rect 111996 114436 112052 114438
rect 112100 114490 112156 114492
rect 112100 114438 112102 114490
rect 112102 114438 112154 114490
rect 112154 114438 112156 114490
rect 112100 114436 112156 114438
rect 112204 114490 112260 114492
rect 112204 114438 112206 114490
rect 112206 114438 112258 114490
rect 112258 114438 112260 114490
rect 112204 114436 112260 114438
rect 111996 112922 112052 112924
rect 111996 112870 111998 112922
rect 111998 112870 112050 112922
rect 112050 112870 112052 112922
rect 111996 112868 112052 112870
rect 112100 112922 112156 112924
rect 112100 112870 112102 112922
rect 112102 112870 112154 112922
rect 112154 112870 112156 112922
rect 112100 112868 112156 112870
rect 112204 112922 112260 112924
rect 112204 112870 112206 112922
rect 112206 112870 112258 112922
rect 112258 112870 112260 112922
rect 112204 112868 112260 112870
rect 111996 111354 112052 111356
rect 111996 111302 111998 111354
rect 111998 111302 112050 111354
rect 112050 111302 112052 111354
rect 111996 111300 112052 111302
rect 112100 111354 112156 111356
rect 112100 111302 112102 111354
rect 112102 111302 112154 111354
rect 112154 111302 112156 111354
rect 112100 111300 112156 111302
rect 112204 111354 112260 111356
rect 112204 111302 112206 111354
rect 112206 111302 112258 111354
rect 112258 111302 112260 111354
rect 112204 111300 112260 111302
rect 111996 109786 112052 109788
rect 111996 109734 111998 109786
rect 111998 109734 112050 109786
rect 112050 109734 112052 109786
rect 111996 109732 112052 109734
rect 112100 109786 112156 109788
rect 112100 109734 112102 109786
rect 112102 109734 112154 109786
rect 112154 109734 112156 109786
rect 112100 109732 112156 109734
rect 112204 109786 112260 109788
rect 112204 109734 112206 109786
rect 112206 109734 112258 109786
rect 112258 109734 112260 109786
rect 112204 109732 112260 109734
rect 111996 108218 112052 108220
rect 111996 108166 111998 108218
rect 111998 108166 112050 108218
rect 112050 108166 112052 108218
rect 111996 108164 112052 108166
rect 112100 108218 112156 108220
rect 112100 108166 112102 108218
rect 112102 108166 112154 108218
rect 112154 108166 112156 108218
rect 112100 108164 112156 108166
rect 112204 108218 112260 108220
rect 112204 108166 112206 108218
rect 112206 108166 112258 108218
rect 112258 108166 112260 108218
rect 112204 108164 112260 108166
rect 111996 106650 112052 106652
rect 111996 106598 111998 106650
rect 111998 106598 112050 106650
rect 112050 106598 112052 106650
rect 111996 106596 112052 106598
rect 112100 106650 112156 106652
rect 112100 106598 112102 106650
rect 112102 106598 112154 106650
rect 112154 106598 112156 106650
rect 112100 106596 112156 106598
rect 112204 106650 112260 106652
rect 112204 106598 112206 106650
rect 112206 106598 112258 106650
rect 112258 106598 112260 106650
rect 112204 106596 112260 106598
rect 111996 105082 112052 105084
rect 111996 105030 111998 105082
rect 111998 105030 112050 105082
rect 112050 105030 112052 105082
rect 111996 105028 112052 105030
rect 112100 105082 112156 105084
rect 112100 105030 112102 105082
rect 112102 105030 112154 105082
rect 112154 105030 112156 105082
rect 112100 105028 112156 105030
rect 112204 105082 112260 105084
rect 112204 105030 112206 105082
rect 112206 105030 112258 105082
rect 112258 105030 112260 105082
rect 112204 105028 112260 105030
rect 111996 103514 112052 103516
rect 111996 103462 111998 103514
rect 111998 103462 112050 103514
rect 112050 103462 112052 103514
rect 111996 103460 112052 103462
rect 112100 103514 112156 103516
rect 112100 103462 112102 103514
rect 112102 103462 112154 103514
rect 112154 103462 112156 103514
rect 112100 103460 112156 103462
rect 112204 103514 112260 103516
rect 112204 103462 112206 103514
rect 112206 103462 112258 103514
rect 112258 103462 112260 103514
rect 112204 103460 112260 103462
rect 111996 101946 112052 101948
rect 111996 101894 111998 101946
rect 111998 101894 112050 101946
rect 112050 101894 112052 101946
rect 111996 101892 112052 101894
rect 112100 101946 112156 101948
rect 112100 101894 112102 101946
rect 112102 101894 112154 101946
rect 112154 101894 112156 101946
rect 112100 101892 112156 101894
rect 112204 101946 112260 101948
rect 112204 101894 112206 101946
rect 112206 101894 112258 101946
rect 112258 101894 112260 101946
rect 112204 101892 112260 101894
rect 111996 100378 112052 100380
rect 111996 100326 111998 100378
rect 111998 100326 112050 100378
rect 112050 100326 112052 100378
rect 111996 100324 112052 100326
rect 112100 100378 112156 100380
rect 112100 100326 112102 100378
rect 112102 100326 112154 100378
rect 112154 100326 112156 100378
rect 112100 100324 112156 100326
rect 112204 100378 112260 100380
rect 112204 100326 112206 100378
rect 112206 100326 112258 100378
rect 112258 100326 112260 100378
rect 112204 100324 112260 100326
rect 111996 98810 112052 98812
rect 111996 98758 111998 98810
rect 111998 98758 112050 98810
rect 112050 98758 112052 98810
rect 111996 98756 112052 98758
rect 112100 98810 112156 98812
rect 112100 98758 112102 98810
rect 112102 98758 112154 98810
rect 112154 98758 112156 98810
rect 112100 98756 112156 98758
rect 112204 98810 112260 98812
rect 112204 98758 112206 98810
rect 112206 98758 112258 98810
rect 112258 98758 112260 98810
rect 112204 98756 112260 98758
rect 111996 97242 112052 97244
rect 111996 97190 111998 97242
rect 111998 97190 112050 97242
rect 112050 97190 112052 97242
rect 111996 97188 112052 97190
rect 112100 97242 112156 97244
rect 112100 97190 112102 97242
rect 112102 97190 112154 97242
rect 112154 97190 112156 97242
rect 112100 97188 112156 97190
rect 112204 97242 112260 97244
rect 112204 97190 112206 97242
rect 112206 97190 112258 97242
rect 112258 97190 112260 97242
rect 112204 97188 112260 97190
rect 111996 95674 112052 95676
rect 111996 95622 111998 95674
rect 111998 95622 112050 95674
rect 112050 95622 112052 95674
rect 111996 95620 112052 95622
rect 112100 95674 112156 95676
rect 112100 95622 112102 95674
rect 112102 95622 112154 95674
rect 112154 95622 112156 95674
rect 112100 95620 112156 95622
rect 112204 95674 112260 95676
rect 112204 95622 112206 95674
rect 112206 95622 112258 95674
rect 112258 95622 112260 95674
rect 112204 95620 112260 95622
rect 111996 94106 112052 94108
rect 111996 94054 111998 94106
rect 111998 94054 112050 94106
rect 112050 94054 112052 94106
rect 111996 94052 112052 94054
rect 112100 94106 112156 94108
rect 112100 94054 112102 94106
rect 112102 94054 112154 94106
rect 112154 94054 112156 94106
rect 112100 94052 112156 94054
rect 112204 94106 112260 94108
rect 112204 94054 112206 94106
rect 112206 94054 112258 94106
rect 112258 94054 112260 94106
rect 112204 94052 112260 94054
rect 111996 92538 112052 92540
rect 111996 92486 111998 92538
rect 111998 92486 112050 92538
rect 112050 92486 112052 92538
rect 111996 92484 112052 92486
rect 112100 92538 112156 92540
rect 112100 92486 112102 92538
rect 112102 92486 112154 92538
rect 112154 92486 112156 92538
rect 112100 92484 112156 92486
rect 112204 92538 112260 92540
rect 112204 92486 112206 92538
rect 112206 92486 112258 92538
rect 112258 92486 112260 92538
rect 112204 92484 112260 92486
rect 111996 90970 112052 90972
rect 111996 90918 111998 90970
rect 111998 90918 112050 90970
rect 112050 90918 112052 90970
rect 111996 90916 112052 90918
rect 112100 90970 112156 90972
rect 112100 90918 112102 90970
rect 112102 90918 112154 90970
rect 112154 90918 112156 90970
rect 112100 90916 112156 90918
rect 112204 90970 112260 90972
rect 112204 90918 112206 90970
rect 112206 90918 112258 90970
rect 112258 90918 112260 90970
rect 112204 90916 112260 90918
rect 111996 89402 112052 89404
rect 111996 89350 111998 89402
rect 111998 89350 112050 89402
rect 112050 89350 112052 89402
rect 111996 89348 112052 89350
rect 112100 89402 112156 89404
rect 112100 89350 112102 89402
rect 112102 89350 112154 89402
rect 112154 89350 112156 89402
rect 112100 89348 112156 89350
rect 112204 89402 112260 89404
rect 112204 89350 112206 89402
rect 112206 89350 112258 89402
rect 112258 89350 112260 89402
rect 112204 89348 112260 89350
rect 111996 87834 112052 87836
rect 111996 87782 111998 87834
rect 111998 87782 112050 87834
rect 112050 87782 112052 87834
rect 111996 87780 112052 87782
rect 112100 87834 112156 87836
rect 112100 87782 112102 87834
rect 112102 87782 112154 87834
rect 112154 87782 112156 87834
rect 112100 87780 112156 87782
rect 112204 87834 112260 87836
rect 112204 87782 112206 87834
rect 112206 87782 112258 87834
rect 112258 87782 112260 87834
rect 112204 87780 112260 87782
rect 111996 86266 112052 86268
rect 111996 86214 111998 86266
rect 111998 86214 112050 86266
rect 112050 86214 112052 86266
rect 111996 86212 112052 86214
rect 112100 86266 112156 86268
rect 112100 86214 112102 86266
rect 112102 86214 112154 86266
rect 112154 86214 112156 86266
rect 112100 86212 112156 86214
rect 112204 86266 112260 86268
rect 112204 86214 112206 86266
rect 112206 86214 112258 86266
rect 112258 86214 112260 86266
rect 112204 86212 112260 86214
rect 111996 84698 112052 84700
rect 111996 84646 111998 84698
rect 111998 84646 112050 84698
rect 112050 84646 112052 84698
rect 111996 84644 112052 84646
rect 112100 84698 112156 84700
rect 112100 84646 112102 84698
rect 112102 84646 112154 84698
rect 112154 84646 112156 84698
rect 112100 84644 112156 84646
rect 112204 84698 112260 84700
rect 112204 84646 112206 84698
rect 112206 84646 112258 84698
rect 112258 84646 112260 84698
rect 112204 84644 112260 84646
rect 111996 83130 112052 83132
rect 111996 83078 111998 83130
rect 111998 83078 112050 83130
rect 112050 83078 112052 83130
rect 111996 83076 112052 83078
rect 112100 83130 112156 83132
rect 112100 83078 112102 83130
rect 112102 83078 112154 83130
rect 112154 83078 112156 83130
rect 112100 83076 112156 83078
rect 112204 83130 112260 83132
rect 112204 83078 112206 83130
rect 112206 83078 112258 83130
rect 112258 83078 112260 83130
rect 112204 83076 112260 83078
rect 111996 81562 112052 81564
rect 111996 81510 111998 81562
rect 111998 81510 112050 81562
rect 112050 81510 112052 81562
rect 111996 81508 112052 81510
rect 112100 81562 112156 81564
rect 112100 81510 112102 81562
rect 112102 81510 112154 81562
rect 112154 81510 112156 81562
rect 112100 81508 112156 81510
rect 112204 81562 112260 81564
rect 112204 81510 112206 81562
rect 112206 81510 112258 81562
rect 112258 81510 112260 81562
rect 112204 81508 112260 81510
rect 111996 79994 112052 79996
rect 111996 79942 111998 79994
rect 111998 79942 112050 79994
rect 112050 79942 112052 79994
rect 111996 79940 112052 79942
rect 112100 79994 112156 79996
rect 112100 79942 112102 79994
rect 112102 79942 112154 79994
rect 112154 79942 112156 79994
rect 112100 79940 112156 79942
rect 112204 79994 112260 79996
rect 112204 79942 112206 79994
rect 112206 79942 112258 79994
rect 112258 79942 112260 79994
rect 112204 79940 112260 79942
rect 111996 78426 112052 78428
rect 111996 78374 111998 78426
rect 111998 78374 112050 78426
rect 112050 78374 112052 78426
rect 111996 78372 112052 78374
rect 112100 78426 112156 78428
rect 112100 78374 112102 78426
rect 112102 78374 112154 78426
rect 112154 78374 112156 78426
rect 112100 78372 112156 78374
rect 112204 78426 112260 78428
rect 112204 78374 112206 78426
rect 112206 78374 112258 78426
rect 112258 78374 112260 78426
rect 112204 78372 112260 78374
rect 111996 76858 112052 76860
rect 111996 76806 111998 76858
rect 111998 76806 112050 76858
rect 112050 76806 112052 76858
rect 111996 76804 112052 76806
rect 112100 76858 112156 76860
rect 112100 76806 112102 76858
rect 112102 76806 112154 76858
rect 112154 76806 112156 76858
rect 112100 76804 112156 76806
rect 112204 76858 112260 76860
rect 112204 76806 112206 76858
rect 112206 76806 112258 76858
rect 112258 76806 112260 76858
rect 112204 76804 112260 76806
rect 111996 75290 112052 75292
rect 111996 75238 111998 75290
rect 111998 75238 112050 75290
rect 112050 75238 112052 75290
rect 111996 75236 112052 75238
rect 112100 75290 112156 75292
rect 112100 75238 112102 75290
rect 112102 75238 112154 75290
rect 112154 75238 112156 75290
rect 112100 75236 112156 75238
rect 112204 75290 112260 75292
rect 112204 75238 112206 75290
rect 112206 75238 112258 75290
rect 112258 75238 112260 75290
rect 112204 75236 112260 75238
rect 111996 73722 112052 73724
rect 111996 73670 111998 73722
rect 111998 73670 112050 73722
rect 112050 73670 112052 73722
rect 111996 73668 112052 73670
rect 112100 73722 112156 73724
rect 112100 73670 112102 73722
rect 112102 73670 112154 73722
rect 112154 73670 112156 73722
rect 112100 73668 112156 73670
rect 112204 73722 112260 73724
rect 112204 73670 112206 73722
rect 112206 73670 112258 73722
rect 112258 73670 112260 73722
rect 112204 73668 112260 73670
rect 111996 72154 112052 72156
rect 111996 72102 111998 72154
rect 111998 72102 112050 72154
rect 112050 72102 112052 72154
rect 111996 72100 112052 72102
rect 112100 72154 112156 72156
rect 112100 72102 112102 72154
rect 112102 72102 112154 72154
rect 112154 72102 112156 72154
rect 112100 72100 112156 72102
rect 112204 72154 112260 72156
rect 112204 72102 112206 72154
rect 112206 72102 112258 72154
rect 112258 72102 112260 72154
rect 112204 72100 112260 72102
rect 111996 70586 112052 70588
rect 111996 70534 111998 70586
rect 111998 70534 112050 70586
rect 112050 70534 112052 70586
rect 111996 70532 112052 70534
rect 112100 70586 112156 70588
rect 112100 70534 112102 70586
rect 112102 70534 112154 70586
rect 112154 70534 112156 70586
rect 112100 70532 112156 70534
rect 112204 70586 112260 70588
rect 112204 70534 112206 70586
rect 112206 70534 112258 70586
rect 112258 70534 112260 70586
rect 112204 70532 112260 70534
rect 111996 69018 112052 69020
rect 111996 68966 111998 69018
rect 111998 68966 112050 69018
rect 112050 68966 112052 69018
rect 111996 68964 112052 68966
rect 112100 69018 112156 69020
rect 112100 68966 112102 69018
rect 112102 68966 112154 69018
rect 112154 68966 112156 69018
rect 112100 68964 112156 68966
rect 112204 69018 112260 69020
rect 112204 68966 112206 69018
rect 112206 68966 112258 69018
rect 112258 68966 112260 69018
rect 112204 68964 112260 68966
rect 111996 67450 112052 67452
rect 111996 67398 111998 67450
rect 111998 67398 112050 67450
rect 112050 67398 112052 67450
rect 111996 67396 112052 67398
rect 112100 67450 112156 67452
rect 112100 67398 112102 67450
rect 112102 67398 112154 67450
rect 112154 67398 112156 67450
rect 112100 67396 112156 67398
rect 112204 67450 112260 67452
rect 112204 67398 112206 67450
rect 112206 67398 112258 67450
rect 112258 67398 112260 67450
rect 112204 67396 112260 67398
rect 111996 65882 112052 65884
rect 111996 65830 111998 65882
rect 111998 65830 112050 65882
rect 112050 65830 112052 65882
rect 111996 65828 112052 65830
rect 112100 65882 112156 65884
rect 112100 65830 112102 65882
rect 112102 65830 112154 65882
rect 112154 65830 112156 65882
rect 112100 65828 112156 65830
rect 112204 65882 112260 65884
rect 112204 65830 112206 65882
rect 112206 65830 112258 65882
rect 112258 65830 112260 65882
rect 112204 65828 112260 65830
rect 107660 64652 107716 64708
rect 108332 64764 108388 64820
rect 111996 64314 112052 64316
rect 111996 64262 111998 64314
rect 111998 64262 112050 64314
rect 112050 64262 112052 64314
rect 111996 64260 112052 64262
rect 112100 64314 112156 64316
rect 112100 64262 112102 64314
rect 112102 64262 112154 64314
rect 112154 64262 112156 64314
rect 112100 64260 112156 64262
rect 112204 64314 112260 64316
rect 112204 64262 112206 64314
rect 112206 64262 112258 64314
rect 112258 64262 112260 64314
rect 112204 64260 112260 64262
rect 108332 63196 108388 63252
rect 111996 62746 112052 62748
rect 111996 62694 111998 62746
rect 111998 62694 112050 62746
rect 112050 62694 112052 62746
rect 111996 62692 112052 62694
rect 112100 62746 112156 62748
rect 112100 62694 112102 62746
rect 112102 62694 112154 62746
rect 112154 62694 112156 62746
rect 112100 62692 112156 62694
rect 112204 62746 112260 62748
rect 112204 62694 112206 62746
rect 112206 62694 112258 62746
rect 112258 62694 112260 62746
rect 112204 62692 112260 62694
rect 111996 61178 112052 61180
rect 111996 61126 111998 61178
rect 111998 61126 112050 61178
rect 112050 61126 112052 61178
rect 111996 61124 112052 61126
rect 112100 61178 112156 61180
rect 112100 61126 112102 61178
rect 112102 61126 112154 61178
rect 112154 61126 112156 61178
rect 112100 61124 112156 61126
rect 112204 61178 112260 61180
rect 112204 61126 112206 61178
rect 112206 61126 112258 61178
rect 112258 61126 112260 61178
rect 112204 61124 112260 61126
rect 106652 60172 106708 60228
rect 111996 59610 112052 59612
rect 111996 59558 111998 59610
rect 111998 59558 112050 59610
rect 112050 59558 112052 59610
rect 111996 59556 112052 59558
rect 112100 59610 112156 59612
rect 112100 59558 112102 59610
rect 112102 59558 112154 59610
rect 112154 59558 112156 59610
rect 112100 59556 112156 59558
rect 112204 59610 112260 59612
rect 112204 59558 112206 59610
rect 112206 59558 112258 59610
rect 112258 59558 112260 59610
rect 112204 59556 112260 59558
rect 108332 59276 108388 59332
rect 108332 58492 108388 58548
rect 104972 55132 105028 55188
rect 110236 58268 110292 58324
rect 103516 37772 103572 37828
rect 104972 53452 105028 53508
rect 108220 52780 108276 52836
rect 108220 46508 108276 46564
rect 108332 47180 108388 47236
rect 104972 5740 105028 5796
rect 103292 4508 103348 4564
rect 104300 4956 104356 5012
rect 100940 4338 100996 4340
rect 100940 4286 100942 4338
rect 100942 4286 100994 4338
rect 100994 4286 100996 4338
rect 100940 4284 100996 4286
rect 103516 4450 103572 4452
rect 103516 4398 103518 4450
rect 103518 4398 103570 4450
rect 103570 4398 103572 4450
rect 103516 4396 103572 4398
rect 100268 3500 100324 3556
rect 100940 3388 100996 3444
rect 101724 3442 101780 3444
rect 101724 3390 101726 3442
rect 101726 3390 101778 3442
rect 101778 3390 101780 3442
rect 101724 3388 101780 3390
rect 102956 3612 103012 3668
rect 102620 3554 102676 3556
rect 102620 3502 102622 3554
rect 102622 3502 102674 3554
rect 102674 3502 102676 3554
rect 102620 3500 102676 3502
rect 104300 4396 104356 4452
rect 104412 3666 104468 3668
rect 104412 3614 104414 3666
rect 104414 3614 104466 3666
rect 104466 3614 104468 3666
rect 104412 3612 104468 3614
rect 111996 58042 112052 58044
rect 111996 57990 111998 58042
rect 111998 57990 112050 58042
rect 112050 57990 112052 58042
rect 111996 57988 112052 57990
rect 112100 58042 112156 58044
rect 112100 57990 112102 58042
rect 112102 57990 112154 58042
rect 112154 57990 112156 58042
rect 112100 57988 112156 57990
rect 112204 58042 112260 58044
rect 112204 57990 112206 58042
rect 112206 57990 112258 58042
rect 112258 57990 112260 58042
rect 112204 57988 112260 57990
rect 111996 56474 112052 56476
rect 111996 56422 111998 56474
rect 111998 56422 112050 56474
rect 112050 56422 112052 56474
rect 111996 56420 112052 56422
rect 112100 56474 112156 56476
rect 112100 56422 112102 56474
rect 112102 56422 112154 56474
rect 112154 56422 112156 56474
rect 112100 56420 112156 56422
rect 112204 56474 112260 56476
rect 112204 56422 112206 56474
rect 112206 56422 112258 56474
rect 112258 56422 112260 56474
rect 112204 56420 112260 56422
rect 111996 54906 112052 54908
rect 111996 54854 111998 54906
rect 111998 54854 112050 54906
rect 112050 54854 112052 54906
rect 111996 54852 112052 54854
rect 112100 54906 112156 54908
rect 112100 54854 112102 54906
rect 112102 54854 112154 54906
rect 112154 54854 112156 54906
rect 112100 54852 112156 54854
rect 112204 54906 112260 54908
rect 112204 54854 112206 54906
rect 112206 54854 112258 54906
rect 112258 54854 112260 54906
rect 112204 54852 112260 54854
rect 111996 53338 112052 53340
rect 111996 53286 111998 53338
rect 111998 53286 112050 53338
rect 112050 53286 112052 53338
rect 111996 53284 112052 53286
rect 112100 53338 112156 53340
rect 112100 53286 112102 53338
rect 112102 53286 112154 53338
rect 112154 53286 112156 53338
rect 112100 53284 112156 53286
rect 112204 53338 112260 53340
rect 112204 53286 112206 53338
rect 112206 53286 112258 53338
rect 112258 53286 112260 53338
rect 112204 53284 112260 53286
rect 111996 51770 112052 51772
rect 111996 51718 111998 51770
rect 111998 51718 112050 51770
rect 112050 51718 112052 51770
rect 111996 51716 112052 51718
rect 112100 51770 112156 51772
rect 112100 51718 112102 51770
rect 112102 51718 112154 51770
rect 112154 51718 112156 51770
rect 112100 51716 112156 51718
rect 112204 51770 112260 51772
rect 112204 51718 112206 51770
rect 112206 51718 112258 51770
rect 112258 51718 112260 51770
rect 112204 51716 112260 51718
rect 111996 50202 112052 50204
rect 111996 50150 111998 50202
rect 111998 50150 112050 50202
rect 112050 50150 112052 50202
rect 111996 50148 112052 50150
rect 112100 50202 112156 50204
rect 112100 50150 112102 50202
rect 112102 50150 112154 50202
rect 112154 50150 112156 50202
rect 112100 50148 112156 50150
rect 112204 50202 112260 50204
rect 112204 50150 112206 50202
rect 112206 50150 112258 50202
rect 112258 50150 112260 50202
rect 112204 50148 112260 50150
rect 111996 48634 112052 48636
rect 111996 48582 111998 48634
rect 111998 48582 112050 48634
rect 112050 48582 112052 48634
rect 111996 48580 112052 48582
rect 112100 48634 112156 48636
rect 112100 48582 112102 48634
rect 112102 48582 112154 48634
rect 112154 48582 112156 48634
rect 112100 48580 112156 48582
rect 112204 48634 112260 48636
rect 112204 48582 112206 48634
rect 112206 48582 112258 48634
rect 112258 48582 112260 48634
rect 112204 48580 112260 48582
rect 111996 47066 112052 47068
rect 111996 47014 111998 47066
rect 111998 47014 112050 47066
rect 112050 47014 112052 47066
rect 111996 47012 112052 47014
rect 112100 47066 112156 47068
rect 112100 47014 112102 47066
rect 112102 47014 112154 47066
rect 112154 47014 112156 47066
rect 112100 47012 112156 47014
rect 112204 47066 112260 47068
rect 112204 47014 112206 47066
rect 112206 47014 112258 47066
rect 112258 47014 112260 47066
rect 112204 47012 112260 47014
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 110236 35196 110292 35252
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 110012 33964 110068 34020
rect 114380 114882 114436 114884
rect 114380 114830 114382 114882
rect 114382 114830 114434 114882
rect 114434 114830 114436 114882
rect 114380 114828 114436 114830
rect 115164 114882 115220 114884
rect 115164 114830 115166 114882
rect 115166 114830 115218 114882
rect 115218 114830 115220 114882
rect 115164 114828 115220 114830
rect 117852 118188 117908 118244
rect 118188 116508 118244 116564
rect 116844 115276 116900 115332
rect 116284 114940 116340 114996
rect 116284 114268 116340 114324
rect 115500 110908 115556 110964
rect 114940 109282 114996 109284
rect 114940 109230 114942 109282
rect 114942 109230 114994 109282
rect 114994 109230 114996 109282
rect 114940 109228 114996 109230
rect 114940 107714 114996 107716
rect 114940 107662 114942 107714
rect 114942 107662 114994 107714
rect 114994 107662 114996 107714
rect 114940 107660 114996 107662
rect 114492 106258 114548 106260
rect 114492 106206 114494 106258
rect 114494 106206 114546 106258
rect 114546 106206 114548 106258
rect 114492 106204 114548 106206
rect 114940 106258 114996 106260
rect 114940 106206 114942 106258
rect 114942 106206 114994 106258
rect 114994 106206 114996 106258
rect 114940 106204 114996 106206
rect 114940 104578 114996 104580
rect 114940 104526 114942 104578
rect 114942 104526 114994 104578
rect 114994 104526 114996 104578
rect 114940 104524 114996 104526
rect 114828 102450 114884 102452
rect 114828 102398 114830 102450
rect 114830 102398 114882 102450
rect 114882 102398 114884 102450
rect 114828 102396 114884 102398
rect 114492 99820 114548 99876
rect 114828 94610 114884 94612
rect 114828 94558 114830 94610
rect 114830 94558 114882 94610
rect 114882 94558 114884 94610
rect 114828 94556 114884 94558
rect 114492 94220 114548 94276
rect 114380 92930 114436 92932
rect 114380 92878 114382 92930
rect 114382 92878 114434 92930
rect 114434 92878 114436 92930
rect 114380 92876 114436 92878
rect 114940 92930 114996 92932
rect 114940 92878 114942 92930
rect 114942 92878 114994 92930
rect 114994 92878 114996 92930
rect 114940 92876 114996 92878
rect 115388 89516 115444 89572
rect 114940 87330 114996 87332
rect 114940 87278 114942 87330
rect 114942 87278 114994 87330
rect 114994 87278 114996 87330
rect 114940 87276 114996 87278
rect 114380 86658 114436 86660
rect 114380 86606 114382 86658
rect 114382 86606 114434 86658
rect 114434 86606 114436 86658
rect 114380 86604 114436 86606
rect 114940 86658 114996 86660
rect 114940 86606 114942 86658
rect 114942 86606 114994 86658
rect 114994 86606 114996 86658
rect 114940 86604 114996 86606
rect 114492 84812 114548 84868
rect 115388 83468 115444 83524
rect 114828 79378 114884 79380
rect 114828 79326 114830 79378
rect 114830 79326 114882 79378
rect 114882 79326 114884 79378
rect 114828 79324 114884 79326
rect 114828 77810 114884 77812
rect 114828 77758 114830 77810
rect 114830 77758 114882 77810
rect 114882 77758 114884 77810
rect 114828 77756 114884 77758
rect 114380 75682 114436 75684
rect 114380 75630 114382 75682
rect 114382 75630 114434 75682
rect 114434 75630 114436 75682
rect 114380 75628 114436 75630
rect 114940 75682 114996 75684
rect 114940 75630 114942 75682
rect 114942 75630 114994 75682
rect 114994 75630 114996 75682
rect 114940 75628 114996 75630
rect 114828 74226 114884 74228
rect 114828 74174 114830 74226
rect 114830 74174 114882 74226
rect 114882 74174 114884 74226
rect 114828 74172 114884 74174
rect 115836 110348 115892 110404
rect 116284 109228 116340 109284
rect 116284 107660 116340 107716
rect 115836 105644 115892 105700
rect 116284 104300 116340 104356
rect 116620 114268 116676 114324
rect 117068 114322 117124 114324
rect 117068 114270 117070 114322
rect 117070 114270 117122 114322
rect 117122 114270 117124 114322
rect 117068 114268 117124 114270
rect 117740 114828 117796 114884
rect 116508 110908 116564 110964
rect 116060 102060 116116 102116
rect 115836 99596 115892 99652
rect 115836 94892 115892 94948
rect 116060 94220 116116 94276
rect 115836 92876 115892 92932
rect 115948 89628 116004 89684
rect 115836 86156 115892 86212
rect 115836 84812 115892 84868
rect 116284 87554 116340 87556
rect 116284 87502 116286 87554
rect 116286 87502 116338 87554
rect 116338 87502 116340 87554
rect 116284 87500 116340 87502
rect 116844 109282 116900 109284
rect 116844 109230 116846 109282
rect 116846 109230 116898 109282
rect 116898 109230 116900 109282
rect 116844 109228 116900 109230
rect 116844 107714 116900 107716
rect 116844 107662 116846 107714
rect 116846 107662 116898 107714
rect 116898 107662 116900 107714
rect 116844 107660 116900 107662
rect 116844 104300 116900 104356
rect 117068 102114 117124 102116
rect 117068 102062 117070 102114
rect 117070 102062 117122 102114
rect 117122 102062 117124 102114
rect 117068 102060 117124 102062
rect 117068 94274 117124 94276
rect 117068 94222 117070 94274
rect 117070 94222 117122 94274
rect 117122 94222 117124 94274
rect 117068 94220 117124 94222
rect 116956 89682 117012 89684
rect 116956 89630 116958 89682
rect 116958 89630 117010 89682
rect 117010 89630 117012 89682
rect 116956 89628 117012 89630
rect 116844 87500 116900 87556
rect 116844 86828 116900 86884
rect 116172 83356 116228 83412
rect 117068 83410 117124 83412
rect 117068 83358 117070 83410
rect 117070 83358 117122 83410
rect 117122 83358 117124 83410
rect 117068 83356 117124 83358
rect 117292 79884 117348 79940
rect 116060 75404 116116 75460
rect 116172 74002 116228 74004
rect 116172 73950 116174 74002
rect 116174 73950 116226 74002
rect 116226 73950 116228 74002
rect 116172 73948 116228 73950
rect 114380 69410 114436 69412
rect 114380 69358 114382 69410
rect 114382 69358 114434 69410
rect 114434 69358 114436 69410
rect 114380 69356 114436 69358
rect 114940 69410 114996 69412
rect 114940 69358 114942 69410
rect 114942 69358 114994 69410
rect 114994 69358 114996 69410
rect 114940 69356 114996 69358
rect 115164 68796 115220 68852
rect 114156 67228 114212 67284
rect 113932 66946 113988 66948
rect 113932 66894 113934 66946
rect 113934 66894 113986 66946
rect 113986 66894 113988 66946
rect 113932 66892 113988 66894
rect 112700 66108 112756 66164
rect 113484 66162 113540 66164
rect 113484 66110 113486 66162
rect 113486 66110 113538 66162
rect 113538 66110 113540 66162
rect 113484 66108 113540 66110
rect 112700 65548 112756 65604
rect 115948 70418 116004 70420
rect 115948 70366 115950 70418
rect 115950 70366 116002 70418
rect 116002 70366 116004 70418
rect 115948 70364 116004 70366
rect 115500 68796 115556 68852
rect 115836 68684 115892 68740
rect 114156 66274 114212 66276
rect 114156 66222 114158 66274
rect 114158 66222 114210 66274
rect 114210 66222 114212 66274
rect 114156 66220 114212 66222
rect 115052 66274 115108 66276
rect 115052 66222 115054 66274
rect 115054 66222 115106 66274
rect 115106 66222 115108 66274
rect 115052 66220 115108 66222
rect 113932 65714 113988 65716
rect 113932 65662 113934 65714
rect 113934 65662 113986 65714
rect 113986 65662 113988 65714
rect 113932 65660 113988 65662
rect 114492 65660 114548 65716
rect 114828 64818 114884 64820
rect 114828 64766 114830 64818
rect 114830 64766 114882 64818
rect 114882 64766 114884 64818
rect 114828 64764 114884 64766
rect 114828 63308 114884 63364
rect 114828 62076 114884 62132
rect 114940 59948 114996 60004
rect 115276 59778 115332 59780
rect 115276 59726 115278 59778
rect 115278 59726 115330 59778
rect 115330 59726 115332 59778
rect 115276 59724 115332 59726
rect 114940 59388 114996 59444
rect 114828 58546 114884 58548
rect 114828 58494 114830 58546
rect 114830 58494 114882 58546
rect 114882 58494 114884 58546
rect 114828 58492 114884 58494
rect 114492 56194 114548 56196
rect 114492 56142 114494 56194
rect 114494 56142 114546 56194
rect 114546 56142 114548 56194
rect 114492 56140 114548 56142
rect 114940 56140 114996 56196
rect 114380 55244 114436 55300
rect 114940 55298 114996 55300
rect 114940 55246 114942 55298
rect 114942 55246 114994 55298
rect 114994 55246 114996 55298
rect 114940 55244 114996 55246
rect 114380 54572 114436 54628
rect 114940 52834 114996 52836
rect 114940 52782 114942 52834
rect 114942 52782 114994 52834
rect 114994 52782 114996 52834
rect 114940 52780 114996 52782
rect 115612 67340 115668 67396
rect 115948 67116 116004 67172
rect 115612 66780 115668 66836
rect 115612 66162 115668 66164
rect 115612 66110 115614 66162
rect 115614 66110 115666 66162
rect 115666 66110 115668 66162
rect 115612 66108 115668 66110
rect 115500 65996 115556 66052
rect 117180 78540 117236 78596
rect 117068 74002 117124 74004
rect 117068 73950 117070 74002
rect 117070 73950 117122 74002
rect 117122 73950 117124 74002
rect 117068 73948 117124 73950
rect 117068 73388 117124 73444
rect 116508 70364 116564 70420
rect 116396 68796 116452 68852
rect 117404 67116 117460 67172
rect 116956 66780 117012 66836
rect 116060 66162 116116 66164
rect 116060 66110 116062 66162
rect 116062 66110 116114 66162
rect 116114 66110 116116 66162
rect 116060 66108 116116 66110
rect 117404 66274 117460 66276
rect 117404 66222 117406 66274
rect 117406 66222 117458 66274
rect 117458 66222 117460 66274
rect 117404 66220 117460 66222
rect 117292 66108 117348 66164
rect 115948 65884 116004 65940
rect 116172 65100 116228 65156
rect 116956 65100 117012 65156
rect 116172 62636 116228 62692
rect 117068 62636 117124 62692
rect 116172 61292 116228 61348
rect 117068 61346 117124 61348
rect 117068 61294 117070 61346
rect 117070 61294 117122 61346
rect 117122 61294 117124 61346
rect 117068 61292 117124 61294
rect 116284 60620 116340 60676
rect 116844 60674 116900 60676
rect 116844 60622 116846 60674
rect 116846 60622 116898 60674
rect 116898 60622 116900 60674
rect 116844 60620 116900 60622
rect 115836 59778 115892 59780
rect 115836 59726 115838 59778
rect 115838 59726 115890 59778
rect 115890 59726 115892 59778
rect 115836 59724 115892 59726
rect 115836 59276 115892 59332
rect 116172 57932 116228 57988
rect 118076 112642 118132 112644
rect 118076 112590 118078 112642
rect 118078 112590 118130 112642
rect 118130 112590 118132 112642
rect 118076 112588 118132 112590
rect 118076 111522 118132 111524
rect 118076 111470 118078 111522
rect 118078 111470 118130 111522
rect 118130 111470 118132 111522
rect 118076 111468 118132 111470
rect 118076 106818 118132 106820
rect 118076 106766 118078 106818
rect 118078 106766 118130 106818
rect 118130 106766 118132 106818
rect 118076 106764 118132 106766
rect 118076 100940 118132 100996
rect 118076 96236 118132 96292
rect 118076 82348 118132 82404
rect 117964 79884 118020 79940
rect 117964 78540 118020 78596
rect 118076 78092 118132 78148
rect 118076 70754 118132 70756
rect 118076 70702 118078 70754
rect 118078 70702 118130 70754
rect 118130 70702 118132 70754
rect 118076 70700 118132 70702
rect 117068 57932 117124 57988
rect 117964 66892 118020 66948
rect 117740 66220 117796 66276
rect 117852 66162 117908 66164
rect 117852 66110 117854 66162
rect 117854 66110 117906 66162
rect 117906 66110 117908 66162
rect 117852 66108 117908 66110
rect 117628 64876 117684 64932
rect 115836 55970 115892 55972
rect 115836 55918 115838 55970
rect 115838 55918 115890 55970
rect 115890 55918 115892 55970
rect 115836 55916 115892 55918
rect 118076 56642 118132 56644
rect 118076 56590 118078 56642
rect 118078 56590 118130 56642
rect 118130 56590 118132 56642
rect 118076 56588 118132 56590
rect 115836 54572 115892 54628
rect 115500 49868 115556 49924
rect 115500 48524 115556 48580
rect 115500 47852 115556 47908
rect 115388 45276 115444 45332
rect 115164 44828 115220 44884
rect 114940 43426 114996 43428
rect 114940 43374 114942 43426
rect 114942 43374 114994 43426
rect 114994 43374 114996 43426
rect 114940 43372 114996 43374
rect 114380 41970 114436 41972
rect 114380 41918 114382 41970
rect 114382 41918 114434 41970
rect 114434 41918 114436 41970
rect 114380 41916 114436 41918
rect 114940 41970 114996 41972
rect 114940 41918 114942 41970
rect 114942 41918 114994 41970
rect 114994 41918 114996 41970
rect 114940 41916 114996 41918
rect 115500 45164 115556 45220
rect 115388 44492 115444 44548
rect 115836 41858 115892 41860
rect 115836 41806 115838 41858
rect 115838 41806 115890 41858
rect 115890 41806 115892 41858
rect 115836 41804 115892 41806
rect 115276 41132 115332 41188
rect 114828 37772 114884 37828
rect 114492 35698 114548 35700
rect 114492 35646 114494 35698
rect 114494 35646 114546 35698
rect 114546 35646 114548 35698
rect 114492 35644 114548 35646
rect 114940 35698 114996 35700
rect 114940 35646 114942 35698
rect 114942 35646 114994 35698
rect 114994 35646 114996 35698
rect 114940 35644 114996 35646
rect 112588 33516 112644 33572
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 112588 32284 112644 32340
rect 112812 35196 112868 35252
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 110012 21532 110068 21588
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 112364 17612 112420 17668
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 112204 14084 112260 14086
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 112364 5852 112420 5908
rect 114604 34018 114660 34020
rect 114604 33966 114606 34018
rect 114606 33966 114658 34018
rect 114658 33966 114660 34018
rect 114604 33964 114660 33966
rect 115164 33964 115220 34020
rect 114940 32674 114996 32676
rect 114940 32622 114942 32674
rect 114942 32622 114994 32674
rect 114994 32622 114996 32674
rect 114940 32620 114996 32622
rect 115500 40460 115556 40516
rect 116284 52556 116340 52612
rect 116844 52556 116900 52612
rect 116956 48802 117012 48804
rect 116956 48750 116958 48802
rect 116958 48750 117010 48802
rect 117010 48750 117012 48802
rect 116956 48748 117012 48750
rect 117292 48748 117348 48804
rect 116508 45330 116564 45332
rect 116508 45278 116510 45330
rect 116510 45278 116562 45330
rect 116562 45278 116564 45330
rect 116508 45276 116564 45278
rect 116284 43148 116340 43204
rect 116844 43148 116900 43204
rect 116060 40124 116116 40180
rect 118076 46508 118132 46564
rect 117404 45276 117460 45332
rect 118300 115164 118356 115220
rect 118188 43708 118244 43764
rect 116284 39676 116340 39732
rect 117068 39730 117124 39732
rect 117068 39678 117070 39730
rect 117070 39678 117122 39730
rect 117122 39678 117124 39730
rect 117068 39676 117124 39678
rect 115612 39228 115668 39284
rect 115500 33628 115556 33684
rect 115388 32284 115444 32340
rect 114380 30210 114436 30212
rect 114380 30158 114382 30210
rect 114382 30158 114434 30210
rect 114434 30158 114436 30210
rect 114380 30156 114436 30158
rect 114940 29932 114996 29988
rect 114380 26290 114436 26292
rect 114380 26238 114382 26290
rect 114382 26238 114434 26290
rect 114434 26238 114436 26290
rect 114380 26236 114436 26238
rect 114940 26290 114996 26292
rect 114940 26238 114942 26290
rect 114942 26238 114994 26290
rect 114994 26238 114996 26290
rect 114940 26236 114996 26238
rect 114716 24444 114772 24500
rect 114492 15426 114548 15428
rect 114492 15374 114494 15426
rect 114494 15374 114546 15426
rect 114546 15374 114548 15426
rect 114492 15372 114548 15374
rect 114492 14530 114548 14532
rect 114492 14478 114494 14530
rect 114494 14478 114546 14530
rect 114546 14478 114548 14530
rect 114492 14476 114548 14478
rect 114492 8258 114548 8260
rect 114492 8206 114494 8258
rect 114494 8206 114546 8258
rect 114546 8206 114548 8258
rect 114492 8204 114548 8206
rect 113148 5906 113204 5908
rect 113148 5854 113150 5906
rect 113150 5854 113202 5906
rect 113202 5854 113204 5906
rect 113148 5852 113204 5854
rect 111356 5010 111412 5012
rect 111356 4958 111358 5010
rect 111358 4958 111410 5010
rect 111410 4958 111412 5010
rect 111356 4956 111412 4958
rect 111916 5010 111972 5012
rect 111916 4958 111918 5010
rect 111918 4958 111970 5010
rect 111970 4958 111972 5010
rect 111916 4956 111972 4958
rect 112252 4898 112308 4900
rect 112252 4846 112254 4898
rect 112254 4846 112306 4898
rect 112306 4846 112308 4898
rect 112252 4844 112308 4846
rect 113148 4844 113204 4900
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112204 4676 112260 4678
rect 112364 4338 112420 4340
rect 112364 4286 112366 4338
rect 112366 4286 112418 4338
rect 112418 4286 112420 4338
rect 112364 4284 112420 4286
rect 111692 4226 111748 4228
rect 111692 4174 111694 4226
rect 111694 4174 111746 4226
rect 111746 4174 111748 4226
rect 111692 4172 111748 4174
rect 108332 3612 108388 3668
rect 111580 3666 111636 3668
rect 111580 3614 111582 3666
rect 111582 3614 111634 3666
rect 111634 3614 111636 3666
rect 111580 3612 111636 3614
rect 112364 3500 112420 3556
rect 110908 3442 110964 3444
rect 110908 3390 110910 3442
rect 110910 3390 110962 3442
rect 110962 3390 110964 3442
rect 110908 3388 110964 3390
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 112588 3442 112644 3444
rect 112588 3390 112590 3442
rect 112590 3390 112642 3442
rect 112642 3390 112644 3442
rect 112588 3388 112644 3390
rect 115500 30380 115556 30436
rect 117292 39228 117348 39284
rect 118076 38668 118132 38724
rect 116172 36370 116228 36372
rect 116172 36318 116174 36370
rect 116174 36318 116226 36370
rect 116226 36318 116228 36370
rect 116172 36316 116228 36318
rect 117068 36316 117124 36372
rect 117068 35756 117124 35812
rect 115836 35084 115892 35140
rect 116060 33964 116116 34020
rect 117180 33964 117236 34020
rect 116620 32674 116676 32676
rect 116620 32622 116622 32674
rect 116622 32622 116674 32674
rect 116674 32622 116676 32674
rect 116620 32620 116676 32622
rect 118076 34018 118132 34020
rect 118076 33966 118078 34018
rect 118078 33966 118130 34018
rect 118130 33966 118132 34018
rect 118076 33964 118132 33966
rect 116396 32338 116452 32340
rect 116396 32286 116398 32338
rect 116398 32286 116450 32338
rect 116450 32286 116452 32338
rect 116396 32284 116452 32286
rect 115500 30210 115556 30212
rect 115500 30158 115502 30210
rect 115502 30158 115554 30210
rect 115554 30158 115556 30210
rect 115500 30156 115556 30158
rect 116284 29986 116340 29988
rect 116284 29934 116286 29986
rect 116286 29934 116338 29986
rect 116338 29934 116340 29986
rect 116284 29932 116340 29934
rect 115500 27020 115556 27076
rect 116172 26908 116228 26964
rect 117404 29932 117460 29988
rect 117068 26962 117124 26964
rect 117068 26910 117070 26962
rect 117070 26910 117122 26962
rect 117122 26910 117124 26962
rect 117068 26908 117124 26910
rect 115836 25676 115892 25732
rect 115500 22316 115556 22372
rect 115164 20972 115220 21028
rect 115500 18956 115556 19012
rect 114940 15372 114996 15428
rect 115836 14924 115892 14980
rect 114940 14530 114996 14532
rect 114940 14478 114942 14530
rect 114942 14478 114994 14530
rect 114994 14478 114996 14530
rect 114940 14476 114996 14478
rect 115836 14252 115892 14308
rect 114940 12066 114996 12068
rect 114940 12014 114942 12066
rect 114942 12014 114994 12066
rect 114994 12014 114996 12066
rect 114940 12012 114996 12014
rect 116284 11788 116340 11844
rect 116844 11788 116900 11844
rect 118076 16994 118132 16996
rect 118076 16942 118078 16994
rect 118078 16942 118130 16994
rect 118130 16942 118132 16994
rect 118076 16940 118132 16942
rect 115500 9548 115556 9604
rect 114940 8258 114996 8260
rect 114940 8206 114942 8258
rect 114942 8206 114994 8258
rect 114994 8206 114996 8258
rect 114940 8204 114996 8206
rect 115836 8204 115892 8260
rect 115500 6860 115556 6916
rect 114828 6802 114884 6804
rect 114828 6750 114830 6802
rect 114830 6750 114882 6802
rect 114882 6750 114884 6802
rect 114828 6748 114884 6750
rect 116172 6188 116228 6244
rect 116732 6188 116788 6244
rect 114940 5964 114996 6020
rect 115500 5740 115556 5796
rect 113820 3500 113876 3556
rect 114268 3388 114324 3444
rect 114940 4396 114996 4452
rect 116284 4956 116340 5012
rect 116172 4844 116228 4900
rect 117292 4956 117348 5012
rect 117068 4898 117124 4900
rect 117068 4846 117070 4898
rect 117070 4846 117122 4898
rect 117122 4846 117124 4898
rect 117068 4844 117124 4846
rect 116844 4732 116900 4788
rect 117292 4508 117348 4564
rect 117404 4732 117460 4788
rect 116284 4450 116340 4452
rect 116284 4398 116286 4450
rect 116286 4398 116338 4450
rect 116338 4398 116340 4450
rect 116284 4396 116340 4398
rect 117068 4284 117124 4340
rect 118860 4508 118916 4564
rect 117852 4396 117908 4452
rect 117628 4172 117684 4228
rect 116508 3442 116564 3444
rect 116508 3390 116510 3442
rect 116510 3390 116562 3442
rect 116562 3390 116564 3442
rect 116508 3388 116564 3390
rect 114492 1484 114548 1540
rect 117852 3500 117908 3556
rect 118076 2156 118132 2212
<< metal3 >>
rect 119200 119560 119800 119784
rect 200 118916 800 119112
rect 200 118888 2044 118916
rect 728 118860 2044 118888
rect 2100 118860 2110 118916
rect 119200 118244 119800 118440
rect 117842 118188 117852 118244
rect 117908 118216 119800 118244
rect 117908 118188 119336 118216
rect 130 117852 140 117908
rect 196 117852 1820 117908
rect 1876 117852 1886 117908
rect 200 117544 800 117768
rect 200 116872 800 117096
rect 84802 116956 84812 117012
rect 84868 116956 86604 117012
rect 86660 116956 86670 117012
rect 119200 116872 119800 117096
rect 4466 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4750 116844
rect 35186 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35470 116844
rect 65906 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66190 116844
rect 96626 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96910 116844
rect 3378 116620 3388 116676
rect 3444 116620 52108 116676
rect 52164 116620 52174 116676
rect 11778 116508 11788 116564
rect 11844 116508 20972 116564
rect 21028 116508 21038 116564
rect 24322 116508 24332 116564
rect 24388 116508 26012 116564
rect 26068 116508 26078 116564
rect 35522 116508 35532 116564
rect 35588 116508 37436 116564
rect 37492 116508 37502 116564
rect 53218 116508 53228 116564
rect 53284 116508 54012 116564
rect 54068 116508 54078 116564
rect 58146 116508 58156 116564
rect 58212 116508 59500 116564
rect 59556 116508 59566 116564
rect 59938 116508 59948 116564
rect 60004 116508 60508 116564
rect 60564 116508 61740 116564
rect 61796 116508 61806 116564
rect 65314 116508 65324 116564
rect 65380 116508 66444 116564
rect 66500 116508 66510 116564
rect 67330 116508 67340 116564
rect 67396 116508 69132 116564
rect 69188 116508 69198 116564
rect 75394 116508 75404 116564
rect 75460 116508 76972 116564
rect 77028 116508 77038 116564
rect 78082 116508 78092 116564
rect 78148 116508 78988 116564
rect 79044 116508 79054 116564
rect 79762 116508 79772 116564
rect 79828 116508 81564 116564
rect 81620 116508 81630 116564
rect 83458 116508 83468 116564
rect 83524 116508 84812 116564
rect 84868 116508 84878 116564
rect 88162 116508 88172 116564
rect 88228 116508 89068 116564
rect 89124 116508 89134 116564
rect 90850 116508 90860 116564
rect 90916 116508 92652 116564
rect 92708 116508 92718 116564
rect 101602 116508 101612 116564
rect 101668 116508 111804 116564
rect 111860 116508 111870 116564
rect 115714 116508 115724 116564
rect 115780 116508 118188 116564
rect 118244 116508 118254 116564
rect 15698 116396 15708 116452
rect 15764 116396 17388 116452
rect 17444 116396 17454 116452
rect 23538 116396 23548 116452
rect 23604 116396 25340 116452
rect 25396 116396 25406 116452
rect 43474 116396 43484 116452
rect 43540 116396 51212 116452
rect 51268 116396 51278 116452
rect 85250 116396 85260 116452
rect 85316 116396 85932 116452
rect 85988 116396 85998 116452
rect 89842 116396 89852 116452
rect 89908 116396 95900 116452
rect 95956 116396 95966 116452
rect 31490 116284 31500 116340
rect 31556 116284 33068 116340
rect 33124 116284 33134 116340
rect 43138 116284 43148 116340
rect 43204 116284 44044 116340
rect 44100 116284 44110 116340
rect 46946 116284 46956 116340
rect 47012 116284 47628 116340
rect 47684 116284 48748 116340
rect 48804 116284 48814 116340
rect 72034 116284 72044 116340
rect 72100 116284 74396 116340
rect 74452 116284 74462 116340
rect 81218 116284 81228 116340
rect 81284 116284 82572 116340
rect 82628 116284 82638 116340
rect 95106 116284 95116 116340
rect 95172 116284 96908 116340
rect 96964 116284 96974 116340
rect 99362 116284 99372 116340
rect 99428 116284 100828 116340
rect 100884 116284 100894 116340
rect 106866 116284 106876 116340
rect 106932 116284 108668 116340
rect 108724 116284 108734 116340
rect 110898 116284 110908 116340
rect 110964 116284 112812 116340
rect 112868 116284 112878 116340
rect 114818 116284 114828 116340
rect 114884 116284 116508 116340
rect 116564 116284 116574 116340
rect 3042 116172 3052 116228
rect 3108 116172 3836 116228
rect 3892 116172 3902 116228
rect 48066 116172 48076 116228
rect 48132 116172 55468 116228
rect 75506 116172 75516 116228
rect 75572 116172 76188 116228
rect 76244 116172 76254 116228
rect 55412 116116 55468 116172
rect 43586 116060 43596 116116
rect 43652 116060 48524 116116
rect 48580 116060 48590 116116
rect 55412 116060 56364 116116
rect 56420 116060 56430 116116
rect 19826 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20110 116060
rect 50546 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50830 116060
rect 81266 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81550 116060
rect 111986 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112270 116060
rect 1922 115948 1932 116004
rect 1988 115948 1998 116004
rect 36306 115948 36316 116004
rect 36372 115948 42140 116004
rect 42196 115948 42206 116004
rect 52098 115948 52108 116004
rect 52164 115948 53116 116004
rect 53172 115948 53182 116004
rect 1932 115892 1988 115948
rect 1932 115836 5740 115892
rect 5796 115836 5806 115892
rect 22754 115836 22764 115892
rect 22820 115836 24108 115892
rect 24164 115836 55468 115892
rect 59266 115836 59276 115892
rect 59332 115836 60060 115892
rect 60116 115836 60126 115892
rect 68786 115836 68796 115892
rect 68852 115836 69580 115892
rect 69636 115836 69646 115892
rect 73378 115836 73388 115892
rect 73444 115836 74172 115892
rect 74228 115836 74238 115892
rect 86146 115836 86156 115892
rect 86212 115836 86940 115892
rect 86996 115836 87006 115892
rect 55412 115780 55468 115836
rect 728 115752 4732 115780
rect 200 115724 4732 115752
rect 4788 115724 4798 115780
rect 46498 115724 46508 115780
rect 46564 115724 47964 115780
rect 48020 115724 48030 115780
rect 55412 115724 62972 115780
rect 63028 115724 63038 115780
rect 76738 115724 76748 115780
rect 76804 115724 77532 115780
rect 77588 115724 77598 115780
rect 78754 115724 78764 115780
rect 78820 115724 78988 115780
rect 79044 115724 79054 115780
rect 81890 115724 81900 115780
rect 81956 115724 83244 115780
rect 83300 115724 83310 115780
rect 108770 115724 108780 115780
rect 108836 115724 110124 115780
rect 110180 115724 110190 115780
rect 110338 115724 110348 115780
rect 110404 115724 111244 115780
rect 111300 115724 111310 115780
rect 200 115528 800 115724
rect 12338 115612 12348 115668
rect 12404 115612 23324 115668
rect 23380 115612 23390 115668
rect 70690 115612 70700 115668
rect 70756 115612 71708 115668
rect 71764 115612 72380 115668
rect 72436 115612 87948 115668
rect 88004 115612 88284 115668
rect 88340 115612 88350 115668
rect 119200 115556 119800 115752
rect 5282 115500 5292 115556
rect 5348 115500 9772 115556
rect 9828 115500 10332 115556
rect 10388 115500 11340 115556
rect 11396 115500 11406 115556
rect 32834 115500 32844 115556
rect 32900 115500 33628 115556
rect 33684 115500 37772 115556
rect 37828 115500 37838 115556
rect 38658 115500 38668 115556
rect 38724 115500 41132 115556
rect 41188 115500 41198 115556
rect 64754 115500 64764 115556
rect 64820 115500 65212 115556
rect 65268 115500 66332 115556
rect 66388 115500 67004 115556
rect 67060 115500 67070 115556
rect 100930 115500 100940 115556
rect 100996 115500 101724 115556
rect 101780 115500 101790 115556
rect 103282 115500 103292 115556
rect 103348 115500 109116 115556
rect 109172 115500 109182 115556
rect 115490 115500 115500 115556
rect 115556 115528 119800 115556
rect 115556 115500 119336 115528
rect 69010 115388 69020 115444
rect 69076 115388 69580 115444
rect 69636 115388 70140 115444
rect 70196 115388 100492 115444
rect 100548 115388 101052 115444
rect 101108 115388 101118 115444
rect 115826 115276 115836 115332
rect 115892 115276 116844 115332
rect 116900 115276 116910 115332
rect 4466 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4750 115276
rect 35186 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35470 115276
rect 65906 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66190 115276
rect 96626 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96910 115276
rect 115490 115164 115500 115220
rect 115556 115164 118300 115220
rect 118356 115164 118366 115220
rect 3154 114940 3164 114996
rect 3220 114940 3612 114996
rect 3668 114940 3836 114996
rect 3892 114940 4396 114996
rect 4452 114940 5292 114996
rect 5348 114940 5358 114996
rect 43586 114940 43596 114996
rect 43652 114940 45388 114996
rect 45444 114940 45454 114996
rect 46386 114940 46396 114996
rect 46452 114940 46956 114996
rect 47012 114940 47022 114996
rect 66994 114940 67004 114996
rect 67060 114940 116284 114996
rect 116340 114940 116350 114996
rect 3042 114828 3052 114884
rect 3108 114828 3724 114884
rect 3780 114828 3790 114884
rect 62962 114828 62972 114884
rect 63028 114828 64428 114884
rect 64484 114828 64494 114884
rect 110786 114828 110796 114884
rect 110852 114828 112588 114884
rect 112644 114828 112654 114884
rect 114370 114828 114380 114884
rect 114436 114828 115164 114884
rect 115220 114828 117740 114884
rect 117796 114828 117806 114884
rect 119200 114856 119800 115080
rect 31892 114716 56924 114772
rect 56980 114716 57484 114772
rect 57540 114716 57550 114772
rect 31892 114660 31948 114716
rect 2370 114604 2380 114660
rect 2436 114604 11900 114660
rect 11956 114604 11966 114660
rect 23314 114604 23324 114660
rect 23380 114604 23772 114660
rect 23828 114604 24668 114660
rect 24724 114604 31948 114660
rect 33954 114604 33964 114660
rect 34020 114604 34860 114660
rect 34916 114604 35532 114660
rect 35588 114604 35598 114660
rect 56466 114604 56476 114660
rect 56532 114604 61292 114660
rect 61348 114604 61358 114660
rect 19826 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20110 114492
rect 50546 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50830 114492
rect 81266 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81550 114492
rect 111986 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112270 114492
rect 200 114184 800 114408
rect 63634 114268 63644 114324
rect 63700 114268 64092 114324
rect 64148 114268 65212 114324
rect 65268 114268 65278 114324
rect 116274 114268 116284 114324
rect 116340 114268 116620 114324
rect 116676 114268 117068 114324
rect 117124 114268 117134 114324
rect 3714 113932 3724 113988
rect 3780 113932 9212 113988
rect 9268 113932 9278 113988
rect 3378 113820 3388 113876
rect 3444 113820 54460 113876
rect 54516 113820 54526 113876
rect 200 113540 800 113736
rect 4466 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4750 113708
rect 35186 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35470 113708
rect 65906 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66190 113708
rect 96626 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96910 113708
rect 200 113512 1820 113540
rect 728 113484 1820 113512
rect 1876 113484 1886 113540
rect 119200 113512 119800 113736
rect 42130 113372 42140 113428
rect 42196 113372 67788 113428
rect 67844 113372 67854 113428
rect 74722 113372 74732 113428
rect 74788 113372 85260 113428
rect 85316 113372 85326 113428
rect 19826 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20110 112924
rect 50546 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50830 112924
rect 81266 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81550 112924
rect 111986 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112270 112924
rect 118066 112588 118076 112644
rect 118132 112588 118142 112644
rect 118076 112420 118132 112588
rect 728 112392 1932 112420
rect 200 112364 1932 112392
rect 1988 112364 1998 112420
rect 118076 112392 119336 112420
rect 118076 112364 119800 112392
rect 200 112168 800 112364
rect 119200 112168 119800 112364
rect 4466 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4750 112140
rect 35186 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35470 112140
rect 65906 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66190 112140
rect 96626 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96910 112140
rect 3266 111804 3276 111860
rect 3332 111804 29372 111860
rect 29428 111804 29438 111860
rect 119200 111524 119800 111720
rect 118066 111468 118076 111524
rect 118132 111496 119800 111524
rect 118132 111468 119336 111496
rect 19826 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20110 111356
rect 50546 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50830 111356
rect 81266 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81550 111356
rect 111986 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112270 111356
rect 728 111048 1708 111076
rect 200 111020 1708 111048
rect 1764 111020 1774 111076
rect 200 110824 800 111020
rect 115490 110908 115500 110964
rect 115556 110908 116508 110964
rect 116564 110908 116574 110964
rect 4466 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4750 110572
rect 35186 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35470 110572
rect 65906 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66190 110572
rect 96626 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96910 110572
rect 115826 110348 115836 110404
rect 115892 110376 119336 110404
rect 115892 110348 119800 110376
rect 119200 110152 119800 110348
rect 19826 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20110 109788
rect 50546 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50830 109788
rect 81266 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81550 109788
rect 111986 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112270 109788
rect 728 109704 1820 109732
rect 200 109676 1820 109704
rect 1876 109676 1886 109732
rect 200 109480 800 109676
rect 93202 109228 93212 109284
rect 93268 109228 114940 109284
rect 114996 109228 115006 109284
rect 116274 109228 116284 109284
rect 116340 109228 116844 109284
rect 116900 109228 116910 109284
rect 116844 109060 116900 109228
rect 116844 109032 119336 109060
rect 200 108808 800 109032
rect 116844 109004 119800 109032
rect 4466 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4750 109004
rect 35186 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35470 109004
rect 65906 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66190 109004
rect 96626 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96910 109004
rect 119200 108808 119800 109004
rect 19826 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20110 108220
rect 50546 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50830 108220
rect 81266 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81550 108220
rect 111986 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112270 108220
rect 728 107688 1820 107716
rect 200 107660 1820 107688
rect 1876 107660 1886 107716
rect 106642 107660 106652 107716
rect 106708 107660 114940 107716
rect 114996 107660 115006 107716
rect 116274 107660 116284 107716
rect 116340 107660 116844 107716
rect 116900 107688 119336 107716
rect 116900 107660 119800 107688
rect 200 107464 800 107660
rect 119200 107464 119800 107660
rect 4466 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4750 107436
rect 35186 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35470 107436
rect 65906 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66190 107436
rect 96626 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96910 107436
rect 119200 106820 119800 107016
rect 118066 106764 118076 106820
rect 118132 106792 119800 106820
rect 118132 106764 119336 106792
rect 19826 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20110 106652
rect 50546 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50830 106652
rect 81266 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81550 106652
rect 111986 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112270 106652
rect 200 106120 800 106344
rect 73938 106204 73948 106260
rect 74004 106204 114492 106260
rect 114548 106204 114940 106260
rect 114996 106204 115006 106260
rect 4466 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4750 105868
rect 35186 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35470 105868
rect 65906 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66190 105868
rect 96626 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96910 105868
rect 45266 105756 45276 105812
rect 45332 105756 46508 105812
rect 46564 105756 46574 105812
rect 200 105448 800 105672
rect 115826 105644 115836 105700
rect 115892 105672 119336 105700
rect 115892 105644 119800 105672
rect 119200 105448 119800 105644
rect 52434 105196 52444 105252
rect 52500 105196 99820 105252
rect 99876 105196 99886 105252
rect 19826 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20110 105084
rect 50546 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50830 105084
rect 81266 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81550 105084
rect 111986 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112270 105084
rect 3042 104524 3052 104580
rect 3108 104524 3612 104580
rect 3668 104524 32732 104580
rect 32788 104524 32798 104580
rect 100034 104524 100044 104580
rect 100100 104524 114940 104580
rect 114996 104524 115006 104580
rect 728 104328 1932 104356
rect 200 104300 1932 104328
rect 1988 104300 1998 104356
rect 116274 104300 116284 104356
rect 116340 104300 116844 104356
rect 116900 104328 119336 104356
rect 116900 104300 119800 104328
rect 200 104104 800 104300
rect 4466 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4750 104300
rect 35186 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35470 104300
rect 65906 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66190 104300
rect 96626 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96910 104300
rect 119200 104104 119800 104300
rect 19826 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20110 103516
rect 50546 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50830 103516
rect 81266 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81550 103516
rect 111986 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112270 103516
rect 728 102984 1932 103012
rect 200 102956 1932 102984
rect 1988 102956 1998 103012
rect 3042 102956 3052 103012
rect 3108 102956 3612 103012
rect 3668 102956 44828 103012
rect 44884 102956 44894 103012
rect 45154 102956 45164 103012
rect 45220 102956 45612 103012
rect 45668 102956 45948 103012
rect 46004 102956 73948 103012
rect 74004 102956 74014 103012
rect 200 102760 800 102956
rect 119200 102760 119800 102984
rect 4466 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4750 102732
rect 35186 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35470 102732
rect 65906 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66190 102732
rect 96626 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96910 102732
rect 3154 102396 3164 102452
rect 3220 102396 22652 102452
rect 22708 102396 22718 102452
rect 56914 102396 56924 102452
rect 56980 102396 114828 102452
rect 114884 102396 114894 102452
rect 119200 102116 119800 102312
rect 116050 102060 116060 102116
rect 116116 102060 117068 102116
rect 117124 102088 119800 102116
rect 117124 102060 119336 102088
rect 19826 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20110 101948
rect 50546 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50830 101948
rect 81266 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81550 101948
rect 111986 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112270 101948
rect 32162 101724 32172 101780
rect 32228 101724 39564 101780
rect 39620 101724 39630 101780
rect 728 101640 2380 101668
rect 200 101612 2380 101640
rect 2436 101612 2446 101668
rect 200 101416 800 101612
rect 4466 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4750 101164
rect 35186 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35470 101164
rect 65906 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66190 101164
rect 96626 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96910 101164
rect 728 100968 1820 100996
rect 200 100940 1820 100968
rect 1876 100940 1886 100996
rect 118066 100940 118076 100996
rect 118132 100968 119336 100996
rect 118132 100940 119800 100968
rect 200 100744 800 100940
rect 119200 100744 119800 100940
rect 19826 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20110 100380
rect 50546 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50830 100380
rect 81266 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81550 100380
rect 111986 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112270 100380
rect 3266 99820 3276 99876
rect 3332 99820 37884 99876
rect 37940 99820 37950 99876
rect 83122 99820 83132 99876
rect 83188 99820 114492 99876
rect 114548 99820 114558 99876
rect 200 99428 800 99624
rect 115826 99596 115836 99652
rect 115892 99624 119336 99652
rect 115892 99596 119800 99624
rect 4466 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4750 99596
rect 35186 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35470 99596
rect 65906 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66190 99596
rect 96626 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96910 99596
rect 200 99400 1820 99428
rect 728 99372 1820 99400
rect 1876 99372 1886 99428
rect 38546 99372 38556 99428
rect 38612 99372 39452 99428
rect 39508 99372 39518 99428
rect 119200 99400 119800 99596
rect 2594 99148 2604 99204
rect 2660 99148 3164 99204
rect 3220 99148 3230 99204
rect 38882 99148 38892 99204
rect 38948 99148 41692 99204
rect 41748 99148 41758 99204
rect 19826 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20110 98812
rect 50546 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50830 98812
rect 81266 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81550 98812
rect 111986 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112270 98812
rect 119200 98728 119800 98952
rect 728 98280 1932 98308
rect 200 98252 1932 98280
rect 1988 98252 1998 98308
rect 200 98056 800 98252
rect 4466 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4750 98028
rect 35186 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35470 98028
rect 65906 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66190 98028
rect 96626 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96910 98028
rect 3266 97692 3276 97748
rect 3332 97692 15932 97748
rect 15988 97692 15998 97748
rect 119200 97384 119800 97608
rect 19826 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20110 97244
rect 50546 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50830 97244
rect 81266 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81550 97244
rect 111986 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112270 97244
rect 728 96936 1708 96964
rect 200 96908 1708 96936
rect 1764 96908 1774 96964
rect 200 96712 800 96908
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 65906 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66190 96460
rect 96626 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96910 96460
rect 200 96040 800 96264
rect 118066 96236 118076 96292
rect 118132 96264 119336 96292
rect 118132 96236 119800 96264
rect 119200 96040 119800 96236
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 50546 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50830 95676
rect 81266 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81550 95676
rect 111986 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112270 95676
rect 728 94920 1932 94948
rect 200 94892 1932 94920
rect 1988 94892 1998 94948
rect 115826 94892 115836 94948
rect 115892 94920 119336 94948
rect 115892 94892 119800 94920
rect 200 94696 800 94892
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 65906 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66190 94892
rect 96626 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96910 94892
rect 119200 94696 119800 94892
rect 88162 94556 88172 94612
rect 88228 94556 114828 94612
rect 114884 94556 114894 94612
rect 61282 94332 61292 94388
rect 61348 94332 71260 94388
rect 71316 94332 71820 94388
rect 71876 94332 71886 94388
rect 72146 94220 72156 94276
rect 72212 94220 114492 94276
rect 114548 94220 114558 94276
rect 116050 94220 116060 94276
rect 116116 94220 117068 94276
rect 117124 94248 119336 94276
rect 117124 94220 119800 94248
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 50546 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50830 94108
rect 81266 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81550 94108
rect 111986 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112270 94108
rect 119200 94024 119800 94220
rect 728 93576 1932 93604
rect 200 93548 1932 93576
rect 1988 93548 1998 93604
rect 3042 93548 3052 93604
rect 3108 93548 3612 93604
rect 3668 93548 48300 93604
rect 48356 93548 48366 93604
rect 48626 93548 48636 93604
rect 48692 93548 49420 93604
rect 49476 93548 61852 93604
rect 61908 93548 67228 93604
rect 200 93352 800 93548
rect 67172 93492 67228 93548
rect 67172 93436 74732 93492
rect 74788 93436 74798 93492
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 65906 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66190 93324
rect 96626 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96910 93324
rect 3266 92988 3276 93044
rect 3332 92988 57932 93044
rect 57988 92988 57998 93044
rect 200 92820 800 92904
rect 98242 92876 98252 92932
rect 98308 92876 114380 92932
rect 114436 92876 114940 92932
rect 114996 92876 115006 92932
rect 115826 92876 115836 92932
rect 115892 92904 119336 92932
rect 115892 92876 119800 92904
rect 200 92764 1932 92820
rect 1988 92764 1998 92820
rect 200 92680 800 92764
rect 119200 92680 119800 92876
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 50546 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50830 92540
rect 81266 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81550 92540
rect 111986 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112270 92540
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 65906 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66190 91756
rect 96626 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96910 91756
rect 200 91336 800 91560
rect 119200 91336 119800 91560
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 50546 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50830 90972
rect 81266 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81550 90972
rect 111986 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112270 90972
rect 119200 90664 119800 90888
rect 728 90216 1932 90244
rect 200 90188 1932 90216
rect 1988 90188 1998 90244
rect 200 89992 800 90188
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 65906 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66190 90188
rect 96626 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96910 90188
rect 5058 89628 5068 89684
rect 5124 89628 55468 89684
rect 115938 89628 115948 89684
rect 116004 89628 116956 89684
rect 117012 89628 117022 89684
rect 55412 89572 55468 89628
rect 55412 89516 58828 89572
rect 58884 89516 59724 89572
rect 59780 89516 60732 89572
rect 60788 89516 60798 89572
rect 115378 89516 115388 89572
rect 115444 89544 119336 89572
rect 115444 89516 119800 89544
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 50546 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50830 89404
rect 81266 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81550 89404
rect 111986 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112270 89404
rect 119200 89320 119800 89516
rect 3042 88956 3052 89012
rect 3108 88956 3500 89012
rect 3556 88956 5068 89012
rect 5124 88956 5134 89012
rect 728 88872 1932 88900
rect 200 88844 1932 88872
rect 1988 88844 1998 88900
rect 200 88648 800 88844
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 65906 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66190 88620
rect 96626 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96910 88620
rect 3266 88284 3276 88340
rect 3332 88284 24332 88340
rect 24388 88284 24398 88340
rect 200 88116 800 88200
rect 200 88060 1932 88116
rect 1988 88060 1998 88116
rect 200 87976 800 88060
rect 119200 87976 119800 88200
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 50546 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50830 87836
rect 81266 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81550 87836
rect 111986 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112270 87836
rect 116274 87500 116284 87556
rect 116340 87500 116844 87556
rect 116900 87500 116910 87556
rect 74722 87276 74732 87332
rect 74788 87276 114940 87332
rect 114996 87276 115006 87332
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 65906 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66190 87052
rect 96626 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96910 87052
rect 200 86632 800 86856
rect 116834 86828 116844 86884
rect 116900 86856 119336 86884
rect 116900 86828 119800 86856
rect 102452 86604 114380 86660
rect 114436 86604 114940 86660
rect 114996 86604 115006 86660
rect 119200 86632 119800 86828
rect 102452 86436 102508 86604
rect 61954 86380 61964 86436
rect 62020 86380 102508 86436
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 50546 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50830 86268
rect 81266 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81550 86268
rect 111986 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112270 86268
rect 115826 86156 115836 86212
rect 115892 86184 119336 86212
rect 115892 86156 119800 86184
rect 119200 85960 119800 86156
rect 728 85512 1820 85540
rect 200 85484 1820 85512
rect 1876 85484 1886 85540
rect 200 85288 800 85484
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 65906 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66190 85484
rect 96626 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96910 85484
rect 76514 84812 76524 84868
rect 76580 84812 114492 84868
rect 114548 84812 114558 84868
rect 115826 84812 115836 84868
rect 115892 84840 119336 84868
rect 115892 84812 119800 84840
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 50546 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50830 84700
rect 81266 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81550 84700
rect 111986 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112270 84700
rect 119200 84616 119800 84812
rect 728 84168 1820 84196
rect 200 84140 1820 84168
rect 1876 84140 1886 84196
rect 200 83944 800 84140
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 65906 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66190 83916
rect 96626 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96910 83916
rect 200 83272 800 83496
rect 115378 83468 115388 83524
rect 115444 83496 119336 83524
rect 115444 83468 119800 83496
rect 116162 83356 116172 83412
rect 116228 83356 117068 83412
rect 117124 83356 117134 83412
rect 119200 83272 119800 83468
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 50546 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50830 83132
rect 81266 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81550 83132
rect 111986 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112270 83132
rect 118066 82348 118076 82404
rect 118132 82348 118142 82404
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 65906 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66190 82348
rect 96626 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96910 82348
rect 118076 82180 118132 82348
rect 728 82152 1932 82180
rect 200 82124 1932 82152
rect 1988 82124 1998 82180
rect 118076 82152 119336 82180
rect 118076 82124 119800 82152
rect 200 81928 800 82124
rect 119200 81928 119800 82124
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 50546 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50830 81564
rect 81266 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81550 81564
rect 111986 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112270 81564
rect 119200 81256 119800 81480
rect 200 80584 800 80808
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 65906 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66190 80780
rect 96626 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96910 80780
rect 728 80136 1932 80164
rect 200 80108 1932 80136
rect 1988 80108 1998 80164
rect 200 79912 800 80108
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 50546 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50830 79996
rect 81266 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81550 79996
rect 111986 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112270 79996
rect 119200 79940 119800 80136
rect 117282 79884 117292 79940
rect 117348 79884 117964 79940
rect 118020 79912 119800 79940
rect 118020 79884 119336 79912
rect 83234 79324 83244 79380
rect 83300 79324 114828 79380
rect 114884 79324 114894 79380
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 65906 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66190 79212
rect 96626 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96910 79212
rect 200 78708 800 78792
rect 200 78652 1932 78708
rect 1988 78652 1998 78708
rect 200 78568 800 78652
rect 119200 78596 119800 78792
rect 3042 78540 3052 78596
rect 3108 78540 3500 78596
rect 3556 78540 5852 78596
rect 5908 78540 5918 78596
rect 117170 78540 117180 78596
rect 117236 78540 117964 78596
rect 118020 78568 119800 78596
rect 118020 78540 119336 78568
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 50546 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50830 78428
rect 81266 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81550 78428
rect 111986 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112270 78428
rect 118066 78092 118076 78148
rect 118132 78120 119336 78148
rect 118132 78092 119800 78120
rect 119200 77896 119800 78092
rect 62178 77756 62188 77812
rect 62244 77756 114828 77812
rect 114884 77756 114894 77812
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 65906 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66190 77644
rect 96626 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96910 77644
rect 200 77224 800 77448
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 81266 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81550 76860
rect 111986 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112270 76860
rect 119200 76552 119800 76776
rect 4386 76188 4396 76244
rect 4452 76188 26012 76244
rect 26068 76188 26078 76244
rect 728 76104 1932 76132
rect 200 76076 1932 76104
rect 1988 76076 1998 76132
rect 200 75880 800 76076
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 96626 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96910 76076
rect 86482 75628 86492 75684
rect 86548 75628 114380 75684
rect 114436 75628 114940 75684
rect 114996 75628 115006 75684
rect 728 75432 1932 75460
rect 200 75404 1932 75432
rect 1988 75404 1998 75460
rect 116050 75404 116060 75460
rect 116116 75432 119336 75460
rect 116116 75404 119800 75432
rect 200 75208 800 75404
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 81266 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81550 75292
rect 111986 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112270 75292
rect 119200 75208 119800 75404
rect 3266 75068 3276 75124
rect 3332 75068 3342 75124
rect 3276 75012 3332 75068
rect 2818 74956 2828 75012
rect 2884 74956 3332 75012
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 96626 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96910 74508
rect 104962 74172 104972 74228
rect 105028 74172 114828 74228
rect 114884 74172 114894 74228
rect 200 73864 800 74088
rect 116162 73948 116172 74004
rect 116228 73948 117068 74004
rect 117124 73948 117134 74004
rect 119200 73864 119800 74088
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 81266 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81550 73724
rect 111986 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112270 73724
rect 117058 73388 117068 73444
rect 117124 73416 119336 73444
rect 117124 73388 119800 73416
rect 119200 73192 119800 73388
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 96626 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96910 72940
rect 200 72520 800 72744
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 81266 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81550 72156
rect 111986 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112270 72156
rect 119200 71848 119800 72072
rect 200 71204 800 71400
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 96626 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96910 71372
rect 200 71176 1820 71204
rect 728 71148 1820 71176
rect 1876 71148 1886 71204
rect 3378 70924 3388 70980
rect 3444 70924 10892 70980
rect 10948 70924 10958 70980
rect 200 70504 800 70728
rect 118066 70700 118076 70756
rect 118132 70728 119336 70756
rect 118132 70700 119800 70728
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 81266 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81550 70588
rect 111986 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112270 70588
rect 119200 70504 119800 70700
rect 2818 70364 2828 70420
rect 2884 70364 3388 70420
rect 3444 70364 3454 70420
rect 115938 70364 115948 70420
rect 116004 70364 116508 70420
rect 116564 70364 116574 70420
rect 16818 69916 16828 69972
rect 16884 69916 36876 69972
rect 36932 69916 36942 69972
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 96626 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96910 69804
rect 7522 69692 7532 69748
rect 7588 69692 17612 69748
rect 17668 69692 17678 69748
rect 200 69300 800 69384
rect 102452 69356 114380 69412
rect 114436 69356 114940 69412
rect 114996 69356 115006 69412
rect 200 69244 1932 69300
rect 1988 69244 1998 69300
rect 200 69160 800 69244
rect 102452 69188 102508 69356
rect 68898 69132 68908 69188
rect 68964 69132 102508 69188
rect 119200 69160 119800 69384
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 81266 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81550 69020
rect 111986 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112270 69020
rect 55906 68796 55916 68852
rect 55972 68796 56476 68852
rect 56532 68796 56542 68852
rect 77074 68796 77084 68852
rect 77140 68796 77868 68852
rect 77924 68796 77934 68852
rect 115154 68796 115164 68852
rect 115220 68796 115500 68852
rect 115556 68796 116396 68852
rect 116452 68796 116462 68852
rect 115826 68684 115836 68740
rect 115892 68712 119336 68740
rect 115892 68684 119800 68712
rect 6738 68460 6748 68516
rect 6804 68460 46060 68516
rect 46116 68460 46844 68516
rect 46900 68460 46910 68516
rect 119200 68488 119800 68684
rect 3042 68348 3052 68404
rect 3108 68348 3612 68404
rect 3668 68348 16156 68404
rect 16212 68348 16222 68404
rect 54450 68236 54460 68292
rect 54516 68236 59276 68292
rect 59332 68236 59342 68292
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 96626 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96910 68236
rect 53218 68124 53228 68180
rect 53284 68124 62188 68180
rect 62244 68124 62254 68180
rect 72370 68124 72380 68180
rect 72436 68124 86268 68180
rect 86324 68124 86334 68180
rect 728 68040 1932 68068
rect 200 68012 1932 68040
rect 1988 68012 1998 68068
rect 15922 68012 15932 68068
rect 15988 68012 53900 68068
rect 53956 68012 53966 68068
rect 67330 68012 67340 68068
rect 67396 68012 83132 68068
rect 83188 68012 83198 68068
rect 83346 68012 83356 68068
rect 83412 68012 91196 68068
rect 91252 68012 91262 68068
rect 200 67816 800 68012
rect 60610 67900 60620 67956
rect 60676 67900 61404 67956
rect 61460 67900 61628 67956
rect 61684 67900 61694 67956
rect 62514 67676 62524 67732
rect 62580 67676 64092 67732
rect 64148 67676 64158 67732
rect 56690 67564 56700 67620
rect 56756 67564 57820 67620
rect 57876 67564 60508 67620
rect 60564 67564 60574 67620
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 81266 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81550 67452
rect 111986 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112270 67452
rect 200 67144 800 67368
rect 115602 67340 115612 67396
rect 115668 67368 119336 67396
rect 115668 67340 119800 67368
rect 82338 67228 82348 67284
rect 82404 67228 114156 67284
rect 114212 67228 114222 67284
rect 72370 67172 72380 67228
rect 72436 67172 72446 67228
rect 49522 67116 49532 67172
rect 49588 67116 50540 67172
rect 50596 67116 50606 67172
rect 54898 67116 54908 67172
rect 54964 67116 55692 67172
rect 55748 67116 56252 67172
rect 56308 67116 56318 67172
rect 58930 67116 58940 67172
rect 58996 67116 63532 67172
rect 63588 67116 63980 67172
rect 64036 67116 64046 67172
rect 64530 67116 64540 67172
rect 64596 67116 64606 67172
rect 72146 67116 72156 67172
rect 72212 67116 72436 67172
rect 115938 67116 115948 67172
rect 116004 67116 117404 67172
rect 117460 67116 117470 67172
rect 119200 67144 119800 67340
rect 64540 67060 64596 67116
rect 48402 67004 48412 67060
rect 48468 67004 49644 67060
rect 49700 67004 49710 67060
rect 51986 67004 51996 67060
rect 52052 67004 52668 67060
rect 52724 67004 55244 67060
rect 55300 67004 57596 67060
rect 57652 67004 59052 67060
rect 59108 67004 60620 67060
rect 60676 67004 61292 67060
rect 61348 67004 62076 67060
rect 62132 67004 62972 67060
rect 63028 67004 65324 67060
rect 65380 67004 65660 67060
rect 65716 67004 65726 67060
rect 72258 67004 72268 67060
rect 72324 67004 73276 67060
rect 73332 67004 73342 67060
rect 47954 66892 47964 66948
rect 48020 66892 50764 66948
rect 50820 66892 50830 66948
rect 55570 66892 55580 66948
rect 55636 66892 56364 66948
rect 56420 66892 56430 66948
rect 74274 66892 74284 66948
rect 74340 66892 74956 66948
rect 75012 66892 77644 66948
rect 77700 66892 78316 66948
rect 78372 66892 80444 66948
rect 80500 66892 81228 66948
rect 81284 66892 113932 66948
rect 113988 66892 117964 66948
rect 118020 66892 118030 66948
rect 50372 66780 70252 66836
rect 70308 66780 72380 66836
rect 72436 66780 74620 66836
rect 74676 66780 74686 66836
rect 115602 66780 115612 66836
rect 115668 66780 116956 66836
rect 117012 66780 117022 66836
rect 50372 66724 50428 66780
rect 46386 66668 46396 66724
rect 46452 66668 50428 66724
rect 50754 66668 50764 66724
rect 50820 66668 51324 66724
rect 51380 66668 62636 66724
rect 62692 66668 62702 66724
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 96626 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96910 66668
rect 32722 66444 32732 66500
rect 32788 66444 44604 66500
rect 44660 66444 44670 66500
rect 47292 66444 49532 66500
rect 49588 66444 49598 66500
rect 54786 66444 54796 66500
rect 54852 66444 56140 66500
rect 56196 66444 56588 66500
rect 56644 66444 56654 66500
rect 60498 66444 60508 66500
rect 60564 66444 70700 66500
rect 70756 66444 71708 66500
rect 71764 66444 71774 66500
rect 73266 66444 73276 66500
rect 73332 66444 74172 66500
rect 74228 66444 83356 66500
rect 83412 66444 83422 66500
rect 47292 66388 47348 66444
rect 3266 66332 3276 66388
rect 3332 66332 32172 66388
rect 32228 66332 32238 66388
rect 36642 66332 36652 66388
rect 36708 66332 47292 66388
rect 47348 66332 47358 66388
rect 48626 66332 48636 66388
rect 48692 66332 49420 66388
rect 49476 66332 49486 66388
rect 55906 66332 55916 66388
rect 55972 66332 59388 66388
rect 59444 66332 59454 66388
rect 78866 66332 78876 66388
rect 78932 66332 79548 66388
rect 79604 66332 80556 66388
rect 80612 66332 80622 66388
rect 31892 66220 53844 66276
rect 54226 66220 54236 66276
rect 54292 66220 57596 66276
rect 57652 66220 57662 66276
rect 57922 66220 57932 66276
rect 57988 66220 58716 66276
rect 58772 66220 58782 66276
rect 74610 66220 74620 66276
rect 74676 66220 75628 66276
rect 75684 66220 77420 66276
rect 77476 66220 78428 66276
rect 78484 66220 78494 66276
rect 78642 66220 78652 66276
rect 78708 66220 82236 66276
rect 82292 66220 82302 66276
rect 114146 66220 114156 66276
rect 114212 66220 115052 66276
rect 115108 66220 115118 66276
rect 117394 66220 117404 66276
rect 117460 66220 117740 66276
rect 117796 66220 117806 66276
rect 31892 66164 31948 66220
rect 12898 66108 12908 66164
rect 12964 66108 31948 66164
rect 51874 66108 51884 66164
rect 51940 66108 52332 66164
rect 52388 66108 52398 66164
rect 53788 66052 53844 66220
rect 54002 66108 54012 66164
rect 54068 66108 55356 66164
rect 55412 66108 55422 66164
rect 67106 66108 67116 66164
rect 67172 66108 77196 66164
rect 77252 66108 78204 66164
rect 78260 66108 78270 66164
rect 112690 66108 112700 66164
rect 112756 66108 113484 66164
rect 113540 66108 115612 66164
rect 115668 66108 115678 66164
rect 116050 66108 116060 66164
rect 116116 66108 117292 66164
rect 117348 66108 117852 66164
rect 117908 66108 117918 66164
rect 78204 66052 78260 66108
rect 200 65828 800 66024
rect 50642 65996 50652 66052
rect 50708 65996 51996 66052
rect 52052 65996 52062 66052
rect 53788 65996 55804 66052
rect 55860 65996 56476 66052
rect 56532 65996 56542 66052
rect 64082 65996 64092 66052
rect 64148 65996 64652 66052
rect 64708 65996 65324 66052
rect 65380 65996 65884 66052
rect 65940 65996 66332 66052
rect 66388 65996 70476 66052
rect 70532 65996 70542 66052
rect 78204 65996 81676 66052
rect 81732 65996 82012 66052
rect 82068 65996 82078 66052
rect 115490 65996 115500 66052
rect 115556 66024 119336 66052
rect 115556 65996 119800 66024
rect 54674 65884 54684 65940
rect 54740 65884 54908 65940
rect 54964 65884 56700 65940
rect 56756 65884 56766 65940
rect 63522 65884 63532 65940
rect 63588 65884 64540 65940
rect 64596 65884 74732 65940
rect 74788 65884 74798 65940
rect 112364 65884 115948 65940
rect 116004 65884 116014 65940
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 81266 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81550 65884
rect 111986 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112270 65884
rect 200 65800 1820 65828
rect 728 65772 1820 65800
rect 1876 65772 1886 65828
rect 62132 65772 67228 65828
rect 62132 65716 62188 65772
rect 55122 65660 55132 65716
rect 55188 65660 56364 65716
rect 56420 65660 62188 65716
rect 67172 65716 67228 65772
rect 112364 65716 112420 65884
rect 119200 65800 119800 65996
rect 67172 65660 112420 65716
rect 113922 65660 113932 65716
rect 113988 65660 114492 65716
rect 114548 65660 114558 65716
rect 45826 65548 45836 65604
rect 45892 65548 46732 65604
rect 46788 65548 46798 65604
rect 47506 65436 47516 65492
rect 47572 65436 48636 65492
rect 48692 65436 49532 65492
rect 49588 65436 49980 65492
rect 50036 65436 50046 65492
rect 53330 65436 53340 65492
rect 53396 65436 53900 65492
rect 53956 65436 54572 65492
rect 54628 65436 54638 65492
rect 57820 65380 57876 65660
rect 58706 65548 58716 65604
rect 58772 65548 62300 65604
rect 62356 65548 62366 65604
rect 63970 65548 63980 65604
rect 64036 65548 64988 65604
rect 65044 65548 65054 65604
rect 65650 65548 65660 65604
rect 65716 65548 66780 65604
rect 66836 65548 66846 65604
rect 70690 65548 70700 65604
rect 70756 65548 72156 65604
rect 72212 65548 72222 65604
rect 78418 65548 78428 65604
rect 78484 65548 112700 65604
rect 112756 65548 112766 65604
rect 61516 65492 61572 65548
rect 61506 65436 61516 65492
rect 61572 65436 61582 65492
rect 62402 65436 62412 65492
rect 62468 65436 62478 65492
rect 62412 65380 62468 65436
rect 55906 65324 55916 65380
rect 55972 65324 57484 65380
rect 57540 65324 57550 65380
rect 57810 65324 57820 65380
rect 57876 65324 57886 65380
rect 60946 65324 60956 65380
rect 61012 65324 62468 65380
rect 63186 65324 63196 65380
rect 63252 65324 63868 65380
rect 63924 65324 63934 65380
rect 74162 65324 74172 65380
rect 74228 65324 75180 65380
rect 75236 65324 75246 65380
rect 48738 65212 48748 65268
rect 48804 65212 65772 65268
rect 65828 65212 65838 65268
rect 119200 65156 119800 65352
rect 36866 65100 36876 65156
rect 36932 65100 54236 65156
rect 54292 65100 54302 65156
rect 56690 65100 56700 65156
rect 56756 65100 57372 65156
rect 57428 65100 58044 65156
rect 58100 65100 58110 65156
rect 116162 65100 116172 65156
rect 116228 65100 116956 65156
rect 117012 65128 119800 65156
rect 117012 65100 119336 65128
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 96626 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96910 65100
rect 46722 64876 46732 64932
rect 46788 64876 47628 64932
rect 47684 64876 47964 64932
rect 48020 64876 48030 64932
rect 70466 64876 70476 64932
rect 70532 64876 117628 64932
rect 117684 64876 117694 64932
rect 46834 64764 46844 64820
rect 46900 64764 50428 64820
rect 57922 64764 57932 64820
rect 57988 64764 60172 64820
rect 60228 64764 60238 64820
rect 62626 64764 62636 64820
rect 62692 64764 67340 64820
rect 67396 64764 68012 64820
rect 68068 64764 68078 64820
rect 108322 64764 108332 64820
rect 108388 64764 114828 64820
rect 114884 64764 114894 64820
rect 200 64456 800 64680
rect 14242 64652 14252 64708
rect 14308 64652 36316 64708
rect 36372 64652 36382 64708
rect 45938 64652 45948 64708
rect 46004 64652 47180 64708
rect 47236 64652 47246 64708
rect 50372 64596 50428 64764
rect 55346 64652 55356 64708
rect 55412 64652 55916 64708
rect 55972 64652 55982 64708
rect 56130 64652 56140 64708
rect 56196 64652 58828 64708
rect 58884 64652 60620 64708
rect 60676 64652 60686 64708
rect 65986 64652 65996 64708
rect 66052 64652 68460 64708
rect 68516 64652 69356 64708
rect 69412 64652 71540 64708
rect 91522 64652 91532 64708
rect 91588 64652 107660 64708
rect 107716 64652 107726 64708
rect 44706 64540 44716 64596
rect 44772 64540 46508 64596
rect 46564 64540 46574 64596
rect 46834 64540 46844 64596
rect 46900 64540 47852 64596
rect 47908 64540 48748 64596
rect 48804 64540 48814 64596
rect 50372 64540 57316 64596
rect 57474 64540 57484 64596
rect 57540 64540 58940 64596
rect 58996 64540 59836 64596
rect 59892 64540 59902 64596
rect 69906 64540 69916 64596
rect 69972 64540 70588 64596
rect 70644 64540 70654 64596
rect 48178 64428 48188 64484
rect 48244 64428 50652 64484
rect 50708 64428 51436 64484
rect 51492 64428 51502 64484
rect 53666 64428 53676 64484
rect 53732 64428 54236 64484
rect 54292 64428 54302 64484
rect 57260 64372 57316 64540
rect 71484 64484 71540 64652
rect 62850 64428 62860 64484
rect 62916 64428 63868 64484
rect 63924 64428 63934 64484
rect 65426 64428 65436 64484
rect 65492 64428 66444 64484
rect 66500 64428 66510 64484
rect 67330 64428 67340 64484
rect 67396 64428 68124 64484
rect 68180 64428 70476 64484
rect 70532 64428 71260 64484
rect 71316 64428 71326 64484
rect 71474 64428 71484 64484
rect 71540 64428 71708 64484
rect 71764 64428 71774 64484
rect 57260 64316 59724 64372
rect 59780 64316 64092 64372
rect 64148 64316 65548 64372
rect 65604 64316 66556 64372
rect 66612 64316 74172 64372
rect 74228 64316 74238 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 81266 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81550 64316
rect 111986 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112270 64316
rect 54002 64204 54012 64260
rect 54068 64204 55244 64260
rect 55300 64204 59500 64260
rect 59556 64204 59566 64260
rect 63074 64204 63084 64260
rect 63140 64204 73948 64260
rect 74004 64204 74014 64260
rect 3378 64092 3388 64148
rect 3444 64092 50428 64148
rect 56802 64092 56812 64148
rect 56868 64092 57820 64148
rect 57876 64092 57886 64148
rect 59826 64092 59836 64148
rect 59892 64092 63868 64148
rect 63924 64092 63934 64148
rect 67666 64092 67676 64148
rect 67732 64092 68572 64148
rect 68628 64092 68638 64148
rect 70690 64092 70700 64148
rect 70756 64092 71148 64148
rect 71204 64092 71214 64148
rect 50372 64036 50428 64092
rect 37762 63980 37772 64036
rect 37828 63980 45836 64036
rect 45892 63980 49644 64036
rect 49700 63980 49710 64036
rect 50372 63980 61180 64036
rect 61236 63980 61246 64036
rect 61954 63980 61964 64036
rect 62020 63980 62636 64036
rect 62692 63980 62702 64036
rect 64866 63980 64876 64036
rect 64932 63980 65660 64036
rect 65716 63980 67116 64036
rect 67172 63980 67182 64036
rect 45602 63868 45612 63924
rect 45668 63868 48636 63924
rect 48692 63868 48702 63924
rect 54338 63868 54348 63924
rect 54404 63868 57596 63924
rect 57652 63868 58268 63924
rect 58324 63868 58334 63924
rect 58482 63868 58492 63924
rect 58548 63868 59836 63924
rect 59892 63868 59902 63924
rect 64194 63868 64204 63924
rect 64260 63868 65324 63924
rect 65380 63868 65390 63924
rect 67554 63868 67564 63924
rect 67620 63868 69468 63924
rect 69524 63868 69534 63924
rect 70466 63868 70476 63924
rect 70532 63868 71148 63924
rect 71204 63868 71214 63924
rect 48402 63756 48412 63812
rect 48468 63756 49532 63812
rect 49588 63756 49598 63812
rect 50372 63700 50428 63812
rect 50484 63756 62188 63812
rect 63746 63756 63756 63812
rect 63812 63756 64764 63812
rect 64820 63756 64830 63812
rect 65538 63756 65548 63812
rect 65604 63756 66220 63812
rect 66276 63756 66286 63812
rect 66658 63756 66668 63812
rect 66724 63756 67452 63812
rect 67508 63756 67518 63812
rect 119200 63784 119800 64008
rect 62132 63700 62188 63756
rect 48178 63644 48188 63700
rect 48244 63644 50204 63700
rect 50260 63644 50428 63700
rect 54338 63644 54348 63700
rect 54404 63644 55244 63700
rect 55300 63644 55310 63700
rect 62132 63644 73388 63700
rect 73444 63644 73454 63700
rect 45714 63532 45724 63588
rect 45780 63532 55356 63588
rect 55412 63532 56140 63588
rect 56196 63532 56364 63588
rect 56420 63532 56430 63588
rect 63970 63532 63980 63588
rect 64036 63532 65548 63588
rect 65604 63532 65614 63588
rect 66322 63532 66332 63588
rect 66388 63532 69020 63588
rect 69076 63532 69086 63588
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 96626 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96910 63532
rect 70130 63420 70140 63476
rect 70196 63420 75852 63476
rect 75908 63420 75918 63476
rect 728 63336 1932 63364
rect 200 63308 1932 63336
rect 1988 63308 1998 63364
rect 20962 63308 20972 63364
rect 21028 63308 53452 63364
rect 53508 63308 53518 63364
rect 57698 63308 57708 63364
rect 57764 63308 73108 63364
rect 73266 63308 73276 63364
rect 73332 63308 114828 63364
rect 114884 63308 114894 63364
rect 200 63112 800 63308
rect 73052 63252 73108 63308
rect 5842 63196 5852 63252
rect 5908 63196 48636 63252
rect 48692 63196 50764 63252
rect 50820 63196 50830 63252
rect 58930 63196 58940 63252
rect 58996 63196 60956 63252
rect 61012 63196 61022 63252
rect 66770 63196 66780 63252
rect 66836 63196 68012 63252
rect 68068 63196 69132 63252
rect 69188 63196 69198 63252
rect 73052 63196 108332 63252
rect 108388 63196 108398 63252
rect 55906 63084 55916 63140
rect 55972 63084 57372 63140
rect 57428 63084 58604 63140
rect 58660 63084 58670 63140
rect 59154 63084 59164 63140
rect 59220 63084 59612 63140
rect 59668 63084 73276 63140
rect 73332 63084 73342 63140
rect 58604 63028 58660 63084
rect 50306 62972 50316 63028
rect 50372 62972 50764 63028
rect 50820 62972 50830 63028
rect 58604 62972 61404 63028
rect 61460 62972 62076 63028
rect 62132 62972 62142 63028
rect 68562 62972 68572 63028
rect 68628 62972 69356 63028
rect 69412 62972 70140 63028
rect 70196 62972 70206 63028
rect 49858 62860 49868 62916
rect 49924 62860 62188 62916
rect 62962 62860 62972 62916
rect 63028 62860 63756 62916
rect 63812 62860 63822 62916
rect 64754 62860 64764 62916
rect 64820 62860 65436 62916
rect 65492 62860 65772 62916
rect 65828 62860 68460 62916
rect 68516 62860 69468 62916
rect 69524 62860 69534 62916
rect 62132 62804 62188 62860
rect 62132 62748 67228 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 200 62580 800 62664
rect 67172 62580 67228 62748
rect 81266 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81550 62748
rect 111986 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112270 62748
rect 116162 62636 116172 62692
rect 116228 62636 117068 62692
rect 117124 62664 119336 62692
rect 117124 62636 119800 62664
rect 200 62524 1820 62580
rect 1876 62524 1886 62580
rect 51314 62524 51324 62580
rect 51380 62524 53564 62580
rect 53620 62524 56252 62580
rect 56308 62524 56318 62580
rect 62514 62524 62524 62580
rect 62580 62524 63084 62580
rect 63140 62524 63150 62580
rect 67172 62524 67340 62580
rect 67396 62524 67406 62580
rect 70018 62524 70028 62580
rect 70084 62524 103292 62580
rect 103348 62524 103358 62580
rect 200 62440 800 62524
rect 48066 62412 48076 62468
rect 48132 62412 49196 62468
rect 49252 62412 49532 62468
rect 49588 62412 49868 62468
rect 49924 62412 50092 62468
rect 50148 62412 50158 62468
rect 54786 62412 54796 62468
rect 54852 62412 56700 62468
rect 56756 62412 56766 62468
rect 58034 62412 58044 62468
rect 58100 62412 58940 62468
rect 58996 62412 60620 62468
rect 60676 62412 67564 62468
rect 67620 62412 67630 62468
rect 73378 62412 73388 62468
rect 73444 62412 74172 62468
rect 74228 62412 74238 62468
rect 119200 62440 119800 62636
rect 22642 62300 22652 62356
rect 22708 62300 52892 62356
rect 52948 62300 54460 62356
rect 54516 62300 54526 62356
rect 55010 62300 55020 62356
rect 55076 62300 55916 62356
rect 55972 62300 55982 62356
rect 61506 62300 61516 62356
rect 61572 62300 61852 62356
rect 61908 62300 61918 62356
rect 63634 62300 63644 62356
rect 63700 62300 65660 62356
rect 65716 62300 65726 62356
rect 71138 62300 71148 62356
rect 71204 62300 71372 62356
rect 71428 62300 71708 62356
rect 71764 62300 71774 62356
rect 72370 62300 72380 62356
rect 72436 62300 73500 62356
rect 73556 62300 73566 62356
rect 73714 62300 73724 62356
rect 73780 62300 74508 62356
rect 74564 62300 74732 62356
rect 74788 62300 98252 62356
rect 98308 62300 98318 62356
rect 48850 62188 48860 62244
rect 48916 62188 51324 62244
rect 51380 62188 51390 62244
rect 53330 62188 53340 62244
rect 53396 62188 55244 62244
rect 55300 62188 55468 62244
rect 55524 62188 55534 62244
rect 69570 62188 69580 62244
rect 69636 62188 70588 62244
rect 70644 62188 70924 62244
rect 70980 62188 70990 62244
rect 47730 62076 47740 62132
rect 47796 62076 48300 62132
rect 48356 62076 49308 62132
rect 49364 62076 49374 62132
rect 50418 62076 50428 62132
rect 50484 62076 51100 62132
rect 51156 62076 51166 62132
rect 55570 62076 55580 62132
rect 55636 62076 73948 62132
rect 73892 62020 73948 62076
rect 78932 62076 114828 62132
rect 114884 62076 114894 62132
rect 78932 62020 78988 62076
rect 48514 61964 48524 62020
rect 48580 61964 56140 62020
rect 56196 61964 56206 62020
rect 73892 61964 78988 62020
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 96626 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96910 61964
rect 67442 61852 67452 61908
rect 67508 61852 70028 61908
rect 70084 61852 70094 61908
rect 70802 61852 70812 61908
rect 70868 61852 72156 61908
rect 72212 61852 72222 61908
rect 53778 61740 53788 61796
rect 53844 61740 54124 61796
rect 54180 61740 54190 61796
rect 60274 61740 60284 61796
rect 60340 61740 98252 61796
rect 98308 61740 98318 61796
rect 3042 61628 3052 61684
rect 3108 61628 3612 61684
rect 3668 61628 6748 61684
rect 6804 61628 6814 61684
rect 50418 61628 50428 61684
rect 50484 61628 51212 61684
rect 51268 61628 52444 61684
rect 52500 61628 52510 61684
rect 59378 61628 59388 61684
rect 59444 61628 59500 61684
rect 59556 61628 59566 61684
rect 61170 61628 61180 61684
rect 61236 61628 67900 61684
rect 67956 61628 68348 61684
rect 68404 61628 68414 61684
rect 70354 61628 70364 61684
rect 70420 61628 71148 61684
rect 71204 61628 72044 61684
rect 72100 61628 72110 61684
rect 74498 61628 74508 61684
rect 74564 61628 84140 61684
rect 84196 61628 84206 61684
rect 66658 61516 66668 61572
rect 66724 61516 67228 61572
rect 67284 61516 81116 61572
rect 81172 61516 83020 61572
rect 83076 61516 83086 61572
rect 58146 61404 58156 61460
rect 58212 61404 83244 61460
rect 83300 61404 83310 61460
rect 728 61320 1932 61348
rect 200 61292 1932 61320
rect 1988 61292 1998 61348
rect 24322 61292 24332 61348
rect 24388 61292 52220 61348
rect 52276 61292 54124 61348
rect 54180 61292 54190 61348
rect 66322 61292 66332 61348
rect 66388 61292 67340 61348
rect 67396 61292 67406 61348
rect 70018 61292 70028 61348
rect 70084 61292 70700 61348
rect 70756 61292 70766 61348
rect 71698 61292 71708 61348
rect 71764 61292 73500 61348
rect 73556 61292 74956 61348
rect 75012 61292 75022 61348
rect 116162 61292 116172 61348
rect 116228 61292 117068 61348
rect 117124 61320 119336 61348
rect 117124 61292 119800 61320
rect 200 61096 800 61292
rect 52658 61180 52668 61236
rect 52724 61180 53676 61236
rect 53732 61180 54348 61236
rect 54404 61180 55020 61236
rect 55076 61180 55086 61236
rect 55794 61180 55804 61236
rect 55860 61180 56364 61236
rect 56420 61180 74172 61236
rect 74228 61180 74238 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 81266 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81550 61180
rect 111986 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112270 61180
rect 51090 61068 51100 61124
rect 51156 61068 62188 61124
rect 67666 61068 67676 61124
rect 67732 61068 68124 61124
rect 68180 61068 68190 61124
rect 119200 61096 119800 61292
rect 62132 61012 62188 61068
rect 52658 60956 52668 61012
rect 52724 60956 53788 61012
rect 53844 60956 53854 61012
rect 55010 60956 55020 61012
rect 55076 60956 56364 61012
rect 56420 60956 56430 61012
rect 62132 60956 68572 61012
rect 68628 60956 69356 61012
rect 69412 60956 70476 61012
rect 70532 60956 70542 61012
rect 71922 60956 71932 61012
rect 71988 60956 72380 61012
rect 72436 60956 72446 61012
rect 73602 60956 73612 61012
rect 73668 60956 74284 61012
rect 74340 60956 74350 61012
rect 5842 60844 5852 60900
rect 5908 60844 58044 60900
rect 58100 60844 58380 60900
rect 58436 60844 58446 60900
rect 58818 60844 58828 60900
rect 58884 60844 59612 60900
rect 59668 60844 61852 60900
rect 61908 60844 61918 60900
rect 62412 60844 68012 60900
rect 68068 60844 68078 60900
rect 62412 60788 62468 60844
rect 46050 60732 46060 60788
rect 46116 60732 47068 60788
rect 47124 60732 47134 60788
rect 50194 60732 50204 60788
rect 50260 60732 50988 60788
rect 51044 60732 51054 60788
rect 53554 60732 53564 60788
rect 53620 60732 55356 60788
rect 55412 60732 55422 60788
rect 56130 60732 56140 60788
rect 56196 60732 58324 60788
rect 58482 60732 58492 60788
rect 58548 60732 59164 60788
rect 59220 60732 59230 60788
rect 59490 60732 59500 60788
rect 59556 60732 61292 60788
rect 61348 60732 61358 60788
rect 61954 60732 61964 60788
rect 62020 60732 62412 60788
rect 62468 60732 62478 60788
rect 64978 60732 64988 60788
rect 65044 60732 65324 60788
rect 65380 60732 65390 60788
rect 58268 60676 58324 60732
rect 67564 60676 67620 60844
rect 69804 60788 69860 60956
rect 70242 60844 70252 60900
rect 70308 60844 70924 60900
rect 70980 60844 71988 60900
rect 71932 60788 71988 60844
rect 69794 60732 69804 60788
rect 69860 60732 69870 60788
rect 71922 60732 71932 60788
rect 71988 60732 71998 60788
rect 50306 60620 50316 60676
rect 50372 60620 51548 60676
rect 51604 60620 55468 60676
rect 55524 60620 55534 60676
rect 56914 60620 56924 60676
rect 56980 60620 57708 60676
rect 57764 60620 57774 60676
rect 58268 60620 59052 60676
rect 59108 60620 59118 60676
rect 64866 60620 64876 60676
rect 64932 60620 65212 60676
rect 65268 60620 66668 60676
rect 66724 60620 66734 60676
rect 67554 60620 67564 60676
rect 67620 60620 67630 60676
rect 72258 60620 72268 60676
rect 72324 60620 73612 60676
rect 73668 60620 73678 60676
rect 116274 60620 116284 60676
rect 116340 60620 116844 60676
rect 116900 60648 119336 60676
rect 116900 60620 119800 60648
rect 52882 60508 52892 60564
rect 52948 60508 54012 60564
rect 54068 60508 54078 60564
rect 55346 60508 55356 60564
rect 55412 60508 58156 60564
rect 58212 60508 58222 60564
rect 58482 60508 58492 60564
rect 58548 60508 58604 60564
rect 58660 60508 58940 60564
rect 58996 60508 60844 60564
rect 60900 60508 60910 60564
rect 63634 60508 63644 60564
rect 63700 60508 65436 60564
rect 65492 60508 65502 60564
rect 65650 60508 65660 60564
rect 65716 60508 67228 60564
rect 67284 60508 67294 60564
rect 68684 60508 69468 60564
rect 69524 60508 69534 60564
rect 68684 60452 68740 60508
rect 52994 60396 53004 60452
rect 53060 60396 53900 60452
rect 53956 60396 55020 60452
rect 55076 60396 58716 60452
rect 58772 60396 64092 60452
rect 64148 60396 64158 60452
rect 66994 60396 67004 60452
rect 67060 60396 67900 60452
rect 67956 60396 67966 60452
rect 68674 60396 68684 60452
rect 68740 60396 68750 60452
rect 119200 60424 119800 60620
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 96626 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96910 60396
rect 55458 60284 55468 60340
rect 55524 60284 62188 60340
rect 66770 60284 66780 60340
rect 66836 60284 78988 60340
rect 62132 60228 62188 60284
rect 78932 60228 78988 60284
rect 3378 60172 3388 60228
rect 3444 60172 5852 60228
rect 5908 60172 5918 60228
rect 37762 60172 37772 60228
rect 37828 60172 50428 60228
rect 57250 60172 57260 60228
rect 57316 60172 59948 60228
rect 60004 60172 60956 60228
rect 61012 60172 61292 60228
rect 61348 60172 61358 60228
rect 62132 60172 69356 60228
rect 69412 60172 70364 60228
rect 70420 60172 70430 60228
rect 78932 60172 106652 60228
rect 106708 60172 106718 60228
rect 50372 60116 50428 60172
rect 45266 60060 45276 60116
rect 45332 60060 47964 60116
rect 48020 60060 49196 60116
rect 49252 60060 49262 60116
rect 50372 60060 63532 60116
rect 63588 60060 63868 60116
rect 63924 60060 64428 60116
rect 64484 60060 64494 60116
rect 200 59892 800 59976
rect 20962 59948 20972 60004
rect 21028 59948 31948 60004
rect 48738 59948 48748 60004
rect 48804 59948 49420 60004
rect 49476 59948 50316 60004
rect 50372 59948 50382 60004
rect 51874 59948 51884 60004
rect 51940 59948 53564 60004
rect 53620 59948 53630 60004
rect 55010 59948 55020 60004
rect 55076 59948 55580 60004
rect 55636 59948 56812 60004
rect 56868 59948 57484 60004
rect 57540 59948 57550 60004
rect 57810 59948 57820 60004
rect 57876 59948 58492 60004
rect 58548 59948 58558 60004
rect 59350 59948 59388 60004
rect 59444 59948 59454 60004
rect 59714 59948 59724 60004
rect 59780 59948 60508 60004
rect 60564 59948 60574 60004
rect 69570 59948 69580 60004
rect 69636 59948 76412 60004
rect 76468 59948 76478 60004
rect 76626 59948 76636 60004
rect 76692 59948 114940 60004
rect 114996 59948 115006 60004
rect 31892 59892 31948 59948
rect 200 59836 1932 59892
rect 1988 59836 1998 59892
rect 31892 59836 46620 59892
rect 46676 59836 47404 59892
rect 47460 59836 48524 59892
rect 48580 59836 48590 59892
rect 50194 59836 50204 59892
rect 50260 59836 50876 59892
rect 50932 59836 51772 59892
rect 51828 59836 51838 59892
rect 52770 59836 52780 59892
rect 52836 59836 55132 59892
rect 55188 59836 55468 59892
rect 55524 59836 56924 59892
rect 56980 59836 56990 59892
rect 200 59752 800 59836
rect 38612 59724 58492 59780
rect 58548 59724 60060 59780
rect 60116 59724 60126 59780
rect 70018 59724 70028 59780
rect 70084 59724 70924 59780
rect 70980 59724 70990 59780
rect 71138 59724 71148 59780
rect 71204 59724 73052 59780
rect 73108 59724 73118 59780
rect 115266 59724 115276 59780
rect 115332 59724 115836 59780
rect 115892 59724 115902 59780
rect 38612 59668 38668 59724
rect 58156 59668 58212 59724
rect 32162 59612 32172 59668
rect 32228 59612 38668 59668
rect 48290 59612 48300 59668
rect 48356 59612 48972 59668
rect 49028 59612 49644 59668
rect 49700 59612 49710 59668
rect 56914 59612 56924 59668
rect 56980 59612 57148 59668
rect 57204 59612 57214 59668
rect 58146 59612 58156 59668
rect 58212 59612 58222 59668
rect 61506 59612 61516 59668
rect 61572 59612 73948 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 50978 59500 50988 59556
rect 51044 59500 51324 59556
rect 51380 59500 51390 59556
rect 60498 59500 60508 59556
rect 60564 59500 62636 59556
rect 62692 59500 62702 59556
rect 68562 59500 68572 59556
rect 68628 59500 68908 59556
rect 68964 59500 69692 59556
rect 69748 59500 71484 59556
rect 71540 59500 71550 59556
rect 73892 59444 73948 59612
rect 81266 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81550 59612
rect 111986 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112270 59612
rect 5842 59388 5852 59444
rect 5908 59388 52332 59444
rect 52388 59388 54908 59444
rect 54964 59388 54974 59444
rect 56242 59388 56252 59444
rect 56308 59388 57036 59444
rect 57092 59388 57820 59444
rect 57876 59388 57886 59444
rect 58454 59388 58492 59444
rect 58548 59388 58558 59444
rect 61842 59388 61852 59444
rect 61908 59388 62860 59444
rect 62916 59388 62926 59444
rect 68338 59388 68348 59444
rect 68404 59388 69356 59444
rect 69412 59388 69422 59444
rect 69906 59388 69916 59444
rect 69972 59388 70588 59444
rect 70644 59388 72044 59444
rect 72100 59388 72110 59444
rect 73892 59388 114940 59444
rect 114996 59388 115006 59444
rect 26002 59276 26012 59332
rect 26068 59276 38668 59332
rect 49298 59276 49308 59332
rect 49364 59276 60116 59332
rect 38612 59108 38668 59276
rect 48738 59164 48748 59220
rect 48804 59164 49756 59220
rect 49812 59164 49822 59220
rect 55234 59164 55244 59220
rect 55300 59164 55916 59220
rect 55972 59164 55982 59220
rect 60060 59108 60116 59276
rect 62132 59276 108332 59332
rect 108388 59276 108398 59332
rect 115826 59276 115836 59332
rect 115892 59304 119336 59332
rect 115892 59276 119800 59304
rect 61170 59164 61180 59220
rect 61236 59164 62076 59220
rect 62132 59164 62188 59276
rect 62738 59164 62748 59220
rect 62804 59164 66780 59220
rect 66836 59164 66846 59220
rect 69458 59164 69468 59220
rect 69524 59164 70812 59220
rect 70868 59164 70878 59220
rect 3266 59052 3276 59108
rect 3332 59052 33516 59108
rect 33572 59052 33582 59108
rect 38612 59052 58716 59108
rect 58772 59052 58782 59108
rect 60060 59052 62188 59108
rect 62962 59052 62972 59108
rect 63028 59052 63532 59108
rect 63588 59052 63598 59108
rect 63970 59052 63980 59108
rect 64036 59052 65548 59108
rect 65604 59052 65614 59108
rect 65874 59052 65884 59108
rect 65940 59052 66668 59108
rect 66724 59052 67116 59108
rect 67172 59052 67182 59108
rect 68450 59052 68460 59108
rect 68516 59052 69188 59108
rect 69346 59052 69356 59108
rect 69412 59052 70028 59108
rect 70084 59052 70094 59108
rect 119200 59080 119800 59276
rect 62132 58996 62188 59052
rect 69132 58996 69188 59052
rect 52770 58940 52780 58996
rect 52836 58940 54684 58996
rect 54740 58940 55804 58996
rect 55860 58940 56924 58996
rect 56980 58940 57596 58996
rect 57652 58940 59892 58996
rect 62132 58940 67676 58996
rect 67732 58940 68572 58996
rect 68628 58940 68638 58996
rect 69132 58940 69580 58996
rect 69636 58940 69916 58996
rect 69972 58940 69982 58996
rect 59836 58884 59892 58940
rect 59602 58828 59612 58884
rect 59668 58828 59678 58884
rect 59836 58828 62860 58884
rect 62916 58828 62926 58884
rect 64754 58828 64764 58884
rect 64820 58828 65324 58884
rect 65380 58828 65390 58884
rect 66994 58828 67004 58884
rect 67060 58828 68460 58884
rect 68516 58828 68526 58884
rect 69122 58828 69132 58884
rect 69188 58828 70028 58884
rect 70084 58828 70364 58884
rect 70420 58828 70430 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 59612 58772 59668 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 96626 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96910 58828
rect 54562 58716 54572 58772
rect 54628 58716 56364 58772
rect 56420 58716 57484 58772
rect 57540 58716 57550 58772
rect 59266 58716 59276 58772
rect 59332 58716 59668 58772
rect 61618 58716 61628 58772
rect 61684 58716 62188 58772
rect 62244 58716 62254 58772
rect 66332 58716 86492 58772
rect 86548 58716 86558 58772
rect 66332 58660 66388 58716
rect 200 58548 800 58632
rect 52210 58604 52220 58660
rect 52276 58604 54460 58660
rect 54516 58604 55356 58660
rect 55412 58604 55422 58660
rect 58594 58604 58604 58660
rect 58660 58604 59388 58660
rect 59444 58604 59948 58660
rect 60004 58604 60014 58660
rect 62514 58604 62524 58660
rect 62580 58604 66388 58660
rect 69794 58604 69804 58660
rect 69860 58604 69870 58660
rect 69804 58548 69860 58604
rect 200 58492 1820 58548
rect 1876 58492 1886 58548
rect 49074 58492 49084 58548
rect 49140 58492 49644 58548
rect 49700 58492 49710 58548
rect 53778 58492 53788 58548
rect 53844 58492 62076 58548
rect 62132 58492 62142 58548
rect 68562 58492 68572 58548
rect 68628 58492 69580 58548
rect 69636 58492 73948 58548
rect 108322 58492 108332 58548
rect 108388 58492 114828 58548
rect 114884 58492 114894 58548
rect 200 58408 800 58492
rect 73892 58436 73948 58492
rect 58258 58380 58268 58436
rect 58324 58380 59164 58436
rect 59220 58380 59230 58436
rect 61394 58380 61404 58436
rect 61460 58380 67228 58436
rect 67284 58380 69244 58436
rect 69300 58380 69310 58436
rect 69458 58380 69468 58436
rect 69524 58380 70924 58436
rect 70980 58380 70990 58436
rect 73892 58380 88508 58436
rect 88564 58380 88574 58436
rect 51986 58268 51996 58324
rect 52052 58268 54460 58324
rect 54516 58268 54526 58324
rect 56018 58268 56028 58324
rect 56084 58268 56700 58324
rect 56756 58268 56766 58324
rect 58706 58268 58716 58324
rect 58772 58268 63756 58324
rect 63812 58268 64876 58324
rect 64932 58268 64942 58324
rect 65538 58268 65548 58324
rect 65604 58268 65772 58324
rect 65828 58268 110236 58324
rect 110292 58268 110302 58324
rect 3490 58156 3500 58212
rect 3556 58156 44492 58212
rect 44548 58156 44558 58212
rect 58370 58156 58380 58212
rect 58436 58156 65884 58212
rect 65940 58156 66220 58212
rect 66276 58156 66286 58212
rect 71250 58156 71260 58212
rect 71316 58156 71708 58212
rect 71764 58156 71774 58212
rect 51314 58044 51324 58100
rect 51380 58044 61404 58100
rect 61460 58044 61470 58100
rect 71362 58044 71372 58100
rect 71428 58044 72044 58100
rect 72100 58044 72110 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 200 57736 800 57960
rect 51324 57876 51380 58044
rect 81266 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81550 58044
rect 111986 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112270 58044
rect 116162 57932 116172 57988
rect 116228 57932 117068 57988
rect 117124 57960 119336 57988
rect 117124 57932 119800 57960
rect 49858 57820 49868 57876
rect 49924 57820 51380 57876
rect 52434 57820 52444 57876
rect 52500 57820 54236 57876
rect 54292 57820 54572 57876
rect 54628 57820 54638 57876
rect 56130 57820 56140 57876
rect 56196 57820 56700 57876
rect 56756 57820 56766 57876
rect 62402 57820 62412 57876
rect 62468 57820 64540 57876
rect 64596 57820 83132 57876
rect 83188 57820 83198 57876
rect 9202 57708 9212 57764
rect 9268 57708 49532 57764
rect 49588 57708 49598 57764
rect 54338 57708 54348 57764
rect 54404 57708 55468 57764
rect 55524 57708 56028 57764
rect 56084 57708 56094 57764
rect 57026 57708 57036 57764
rect 57092 57708 57372 57764
rect 57428 57708 60620 57764
rect 60676 57708 61964 57764
rect 62020 57708 62030 57764
rect 119200 57736 119800 57932
rect 36306 57596 36316 57652
rect 36372 57596 51996 57652
rect 52052 57596 52062 57652
rect 57810 57596 57820 57652
rect 57876 57596 59276 57652
rect 59332 57596 59342 57652
rect 65762 57596 65772 57652
rect 65828 57596 66332 57652
rect 66388 57596 66556 57652
rect 66612 57596 66622 57652
rect 48738 57484 48748 57540
rect 48804 57484 49868 57540
rect 49924 57484 49934 57540
rect 50530 57484 50540 57540
rect 50596 57484 50988 57540
rect 51044 57484 51212 57540
rect 51268 57484 52668 57540
rect 52724 57484 52734 57540
rect 55346 57484 55356 57540
rect 55412 57484 57036 57540
rect 57092 57484 59500 57540
rect 59556 57484 59566 57540
rect 60498 57484 60508 57540
rect 60564 57484 60844 57540
rect 60900 57484 61628 57540
rect 61684 57484 61852 57540
rect 61908 57484 61918 57540
rect 64642 57484 64652 57540
rect 64708 57484 65436 57540
rect 65492 57484 89852 57540
rect 89908 57484 89918 57540
rect 26002 57372 26012 57428
rect 26068 57372 54684 57428
rect 54740 57372 58380 57428
rect 58436 57372 58446 57428
rect 44594 57260 44604 57316
rect 44660 57260 52444 57316
rect 52500 57260 52510 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 96626 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96910 57260
rect 51202 57148 51212 57204
rect 51268 57148 51436 57204
rect 51492 57148 52892 57204
rect 52948 57148 55580 57204
rect 55636 57148 57820 57204
rect 57876 57148 57886 57204
rect 65538 57148 65548 57204
rect 65604 57148 65614 57204
rect 65548 57092 65604 57148
rect 63522 57036 63532 57092
rect 63588 57036 65324 57092
rect 65380 57036 65390 57092
rect 65548 57036 66668 57092
rect 66724 57036 66734 57092
rect 70578 57036 70588 57092
rect 70644 57036 71260 57092
rect 71316 57036 71596 57092
rect 71652 57036 73052 57092
rect 73108 57036 73118 57092
rect 73052 56980 73108 57036
rect 55906 56924 55916 56980
rect 55972 56924 56700 56980
rect 56756 56924 57260 56980
rect 57316 56924 57326 56980
rect 58146 56924 58156 56980
rect 58212 56924 58940 56980
rect 58996 56924 59006 56980
rect 59266 56924 59276 56980
rect 59332 56924 59836 56980
rect 59892 56924 61404 56980
rect 61460 56924 62300 56980
rect 62356 56924 62366 56980
rect 62626 56924 62636 56980
rect 62692 56924 63308 56980
rect 63364 56924 63374 56980
rect 63970 56924 63980 56980
rect 64036 56924 64988 56980
rect 65044 56924 65054 56980
rect 65538 56924 65548 56980
rect 65604 56924 66444 56980
rect 66500 56924 66510 56980
rect 69570 56924 69580 56980
rect 69636 56924 70924 56980
rect 70980 56924 70990 56980
rect 73052 56924 80108 56980
rect 80164 56924 80174 56980
rect 17602 56812 17612 56868
rect 17668 56812 47404 56868
rect 47460 56812 50428 56868
rect 50484 56812 50494 56868
rect 52658 56812 52668 56868
rect 52724 56812 53564 56868
rect 53620 56812 53900 56868
rect 53956 56812 53966 56868
rect 60386 56812 60396 56868
rect 60452 56812 62804 56868
rect 64306 56812 64316 56868
rect 64372 56812 65100 56868
rect 65156 56812 66892 56868
rect 66948 56812 66958 56868
rect 67890 56812 67900 56868
rect 67956 56812 72492 56868
rect 72548 56812 72558 56868
rect 62748 56756 62804 56812
rect 67900 56756 67956 56812
rect 22642 56700 22652 56756
rect 22708 56700 62524 56756
rect 62580 56700 62590 56756
rect 62748 56700 67004 56756
rect 67060 56700 67956 56756
rect 728 56616 1932 56644
rect 200 56588 1932 56616
rect 1988 56588 1998 56644
rect 3042 56588 3052 56644
rect 3108 56588 3500 56644
rect 3556 56588 44940 56644
rect 44996 56588 45006 56644
rect 49970 56588 49980 56644
rect 50036 56588 50876 56644
rect 50932 56588 50942 56644
rect 51538 56588 51548 56644
rect 51604 56588 52220 56644
rect 52276 56588 53340 56644
rect 53396 56588 53406 56644
rect 60050 56588 60060 56644
rect 60116 56588 60732 56644
rect 60788 56588 66332 56644
rect 66388 56588 66398 56644
rect 66658 56588 66668 56644
rect 66724 56588 67452 56644
rect 67508 56588 67518 56644
rect 118066 56588 118076 56644
rect 118132 56616 119336 56644
rect 118132 56588 119800 56616
rect 200 56392 800 56588
rect 62290 56476 62300 56532
rect 62356 56476 63532 56532
rect 63588 56476 64316 56532
rect 64372 56476 64382 56532
rect 65538 56476 65548 56532
rect 65604 56476 67788 56532
rect 67844 56476 68572 56532
rect 68628 56476 69132 56532
rect 69188 56476 69198 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 111986 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112270 56476
rect 36194 56364 36204 56420
rect 36260 56364 48412 56420
rect 48468 56364 49644 56420
rect 49700 56364 49710 56420
rect 53890 56364 53900 56420
rect 53956 56364 55356 56420
rect 55412 56364 78652 56420
rect 78708 56364 78718 56420
rect 119200 56392 119800 56588
rect 44482 56252 44492 56308
rect 44548 56252 51156 56308
rect 52322 56252 52332 56308
rect 52388 56252 56140 56308
rect 56196 56252 56700 56308
rect 56756 56252 57372 56308
rect 57428 56252 57438 56308
rect 62402 56252 62412 56308
rect 62468 56252 64092 56308
rect 64148 56252 64158 56308
rect 68562 56252 68572 56308
rect 68628 56252 69692 56308
rect 69748 56252 69758 56308
rect 70130 56252 70140 56308
rect 70196 56252 70700 56308
rect 70756 56252 71148 56308
rect 71204 56252 71932 56308
rect 71988 56252 71998 56308
rect 78932 56252 79772 56308
rect 79828 56252 79838 56308
rect 51100 56196 51156 56252
rect 78932 56196 78988 56252
rect 46162 56140 46172 56196
rect 46228 56140 47068 56196
rect 47124 56140 47134 56196
rect 48626 56140 48636 56196
rect 48692 56140 50932 56196
rect 51090 56140 51100 56196
rect 51156 56140 54460 56196
rect 54516 56140 54526 56196
rect 63746 56140 63756 56196
rect 63812 56140 64204 56196
rect 64260 56140 78988 56196
rect 80322 56140 80332 56196
rect 80388 56140 114492 56196
rect 114548 56140 114940 56196
rect 114996 56140 115006 56196
rect 50876 56084 50932 56140
rect 46946 56028 46956 56084
rect 47012 56028 47852 56084
rect 47908 56028 48524 56084
rect 48580 56028 48590 56084
rect 48850 56028 48860 56084
rect 48916 56028 50204 56084
rect 50260 56028 50652 56084
rect 50708 56028 50718 56084
rect 50876 56028 52332 56084
rect 52388 56028 52398 56084
rect 53778 56028 53788 56084
rect 53844 56028 54908 56084
rect 54964 56028 54974 56084
rect 57586 56028 57596 56084
rect 57652 56028 59500 56084
rect 59556 56028 59566 56084
rect 60162 56028 60172 56084
rect 60228 56028 60844 56084
rect 60900 56028 60910 56084
rect 68898 56028 68908 56084
rect 68964 56028 71484 56084
rect 71540 56028 71550 56084
rect 33506 55916 33516 55972
rect 33572 55916 45612 55972
rect 45668 55916 48300 55972
rect 48356 55916 51996 55972
rect 52052 55916 52062 55972
rect 53666 55916 53676 55972
rect 53732 55916 56364 55972
rect 56420 55916 56430 55972
rect 62850 55916 62860 55972
rect 62916 55916 63756 55972
rect 63812 55916 64540 55972
rect 64596 55916 64606 55972
rect 65090 55916 65100 55972
rect 65156 55916 65772 55972
rect 65828 55916 65838 55972
rect 68450 55916 68460 55972
rect 68516 55916 71036 55972
rect 71092 55916 71102 55972
rect 71922 55916 71932 55972
rect 71988 55916 72604 55972
rect 72660 55916 72670 55972
rect 115826 55916 115836 55972
rect 115892 55944 119336 55972
rect 115892 55916 119800 55944
rect 41682 55804 41692 55860
rect 41748 55804 50540 55860
rect 50596 55804 50606 55860
rect 50978 55804 50988 55860
rect 51044 55804 51548 55860
rect 51604 55804 51614 55860
rect 52882 55804 52892 55860
rect 52948 55804 55804 55860
rect 55860 55804 55870 55860
rect 56018 55804 56028 55860
rect 56084 55804 59164 55860
rect 59220 55804 59230 55860
rect 67778 55804 67788 55860
rect 67844 55804 68348 55860
rect 68404 55804 93212 55860
rect 93268 55804 93278 55860
rect 47954 55692 47964 55748
rect 48020 55692 49868 55748
rect 49924 55692 51100 55748
rect 51156 55692 51166 55748
rect 51426 55692 51436 55748
rect 51492 55692 53788 55748
rect 53844 55692 60172 55748
rect 60228 55692 60238 55748
rect 66546 55692 66556 55748
rect 66612 55692 67340 55748
rect 67396 55692 88172 55748
rect 88228 55692 88238 55748
rect 119200 55720 119800 55916
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 50278 55580 50316 55636
rect 50372 55580 50382 55636
rect 50642 55580 50652 55636
rect 50708 55580 53452 55636
rect 53508 55580 53518 55636
rect 54674 55580 54684 55636
rect 54740 55580 58940 55636
rect 58996 55580 59006 55636
rect 64866 55580 64876 55636
rect 64932 55580 65548 55636
rect 65604 55580 65614 55636
rect 48290 55468 48300 55524
rect 48356 55468 48636 55524
rect 48692 55468 48702 55524
rect 49186 55468 49196 55524
rect 49252 55468 49644 55524
rect 49700 55468 49710 55524
rect 50082 55468 50092 55524
rect 50148 55468 51884 55524
rect 51940 55468 51950 55524
rect 53106 55468 53116 55524
rect 53172 55468 55132 55524
rect 55188 55468 55198 55524
rect 63970 55468 63980 55524
rect 64036 55468 64652 55524
rect 64708 55468 69356 55524
rect 69412 55468 69422 55524
rect 71474 55468 71484 55524
rect 71540 55468 103516 55524
rect 103572 55468 103582 55524
rect 40002 55356 40012 55412
rect 40068 55356 40908 55412
rect 40964 55356 40974 55412
rect 50372 55356 50820 55412
rect 51986 55356 51996 55412
rect 52052 55356 52332 55412
rect 52388 55356 52398 55412
rect 52546 55356 52556 55412
rect 52612 55356 54124 55412
rect 54180 55356 54190 55412
rect 59378 55356 59388 55412
rect 59444 55356 62076 55412
rect 62132 55356 63644 55412
rect 63700 55356 63710 55412
rect 65986 55356 65996 55412
rect 66052 55356 66668 55412
rect 66724 55356 66734 55412
rect 68114 55356 68124 55412
rect 68180 55356 69692 55412
rect 69748 55356 71708 55412
rect 71764 55356 71774 55412
rect 50372 55300 50428 55356
rect 50764 55300 50820 55356
rect 65996 55300 66052 55356
rect 200 55048 800 55272
rect 40786 55244 40796 55300
rect 40852 55244 48972 55300
rect 49028 55244 49196 55300
rect 49252 55244 50428 55300
rect 50530 55244 50540 55300
rect 50596 55244 50606 55300
rect 50764 55244 53676 55300
rect 53732 55244 53742 55300
rect 56354 55244 56364 55300
rect 56420 55244 59164 55300
rect 59220 55244 59230 55300
rect 61730 55244 61740 55300
rect 61796 55244 62300 55300
rect 62356 55244 62366 55300
rect 62850 55244 62860 55300
rect 62916 55244 66052 55300
rect 68898 55244 68908 55300
rect 68964 55244 70364 55300
rect 70420 55244 70430 55300
rect 70578 55244 70588 55300
rect 70644 55244 71484 55300
rect 71540 55244 101836 55300
rect 101892 55244 101902 55300
rect 114370 55244 114380 55300
rect 114436 55244 114940 55300
rect 114996 55244 115006 55300
rect 50540 55188 50596 55244
rect 70364 55188 70420 55244
rect 50540 55132 53900 55188
rect 53956 55132 62748 55188
rect 62804 55132 62814 55188
rect 62962 55132 62972 55188
rect 63028 55132 65100 55188
rect 65156 55132 65166 55188
rect 68674 55132 68684 55188
rect 68740 55132 69580 55188
rect 69636 55132 69646 55188
rect 70364 55132 71036 55188
rect 71092 55132 71102 55188
rect 73892 55132 104972 55188
rect 105028 55132 105038 55188
rect 73892 55076 73948 55132
rect 24322 55020 24332 55076
rect 24388 55020 39676 55076
rect 39732 55020 40684 55076
rect 40740 55020 40750 55076
rect 42242 55020 42252 55076
rect 42308 55020 43372 55076
rect 43428 55020 48188 55076
rect 48244 55020 50204 55076
rect 50260 55020 50270 55076
rect 51202 55020 51212 55076
rect 51268 55020 52108 55076
rect 52164 55020 52174 55076
rect 52434 55020 52444 55076
rect 52500 55020 57484 55076
rect 57540 55020 57932 55076
rect 57988 55020 57998 55076
rect 58146 55020 58156 55076
rect 58212 55020 58604 55076
rect 58660 55020 59500 55076
rect 59556 55020 59566 55076
rect 62290 55020 62300 55076
rect 62356 55020 63644 55076
rect 63700 55020 63710 55076
rect 69458 55020 69468 55076
rect 69524 55020 71932 55076
rect 71988 55020 73948 55076
rect 47842 54908 47852 54964
rect 47908 54908 49308 54964
rect 49364 54908 49756 54964
rect 49812 54908 49822 54964
rect 50978 54908 50988 54964
rect 51044 54908 51082 54964
rect 51202 54908 51212 54964
rect 51268 54908 51660 54964
rect 51716 54908 51726 54964
rect 55906 54908 55916 54964
rect 55972 54908 58268 54964
rect 58324 54908 58828 54964
rect 58884 54908 58894 54964
rect 60620 54908 62860 54964
rect 62916 54908 62926 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 60620 54852 60676 54908
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 111986 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112270 54908
rect 46498 54796 46508 54852
rect 46564 54796 48188 54852
rect 48244 54796 49084 54852
rect 49140 54796 49532 54852
rect 49588 54796 49598 54852
rect 51762 54796 51772 54852
rect 51828 54796 51866 54852
rect 55122 54796 55132 54852
rect 55188 54796 58492 54852
rect 58548 54796 60620 54852
rect 60676 54796 60686 54852
rect 62738 54796 62748 54852
rect 62804 54796 68012 54852
rect 68068 54796 68460 54852
rect 68516 54796 68526 54852
rect 44930 54684 44940 54740
rect 44996 54684 45724 54740
rect 45780 54684 47292 54740
rect 47348 54684 47358 54740
rect 48850 54684 48860 54740
rect 48916 54684 51548 54740
rect 51604 54684 51614 54740
rect 52210 54684 52220 54740
rect 52276 54684 53004 54740
rect 53060 54684 53070 54740
rect 56690 54684 56700 54740
rect 56756 54684 57820 54740
rect 57876 54684 57886 54740
rect 63858 54684 63868 54740
rect 63924 54684 64428 54740
rect 64484 54684 64494 54740
rect 66322 54684 66332 54740
rect 66388 54684 92988 54740
rect 93044 54684 93054 54740
rect 728 54600 1820 54628
rect 200 54572 1820 54600
rect 1876 54572 1886 54628
rect 40898 54572 40908 54628
rect 40964 54572 41580 54628
rect 41636 54572 41646 54628
rect 45724 54572 46172 54628
rect 46228 54572 46508 54628
rect 46564 54572 46574 54628
rect 49634 54572 49644 54628
rect 49700 54572 62188 54628
rect 63186 54572 63196 54628
rect 63252 54572 66556 54628
rect 66612 54572 66622 54628
rect 66994 54572 67004 54628
rect 67060 54572 68796 54628
rect 68852 54572 76636 54628
rect 76692 54572 76702 54628
rect 89954 54572 89964 54628
rect 90020 54572 114380 54628
rect 114436 54572 114446 54628
rect 115826 54572 115836 54628
rect 115892 54600 119336 54628
rect 115892 54572 119800 54600
rect 200 54376 800 54572
rect 45724 54516 45780 54572
rect 62132 54516 62188 54572
rect 45714 54460 45724 54516
rect 45780 54460 45790 54516
rect 47394 54460 47404 54516
rect 47460 54460 48636 54516
rect 48692 54460 49868 54516
rect 49924 54460 49934 54516
rect 50194 54460 50204 54516
rect 50260 54460 50316 54516
rect 50372 54460 50382 54516
rect 51090 54460 51100 54516
rect 51156 54460 51212 54516
rect 51268 54460 54572 54516
rect 54628 54460 55692 54516
rect 55748 54460 55758 54516
rect 56466 54460 56476 54516
rect 56532 54460 56924 54516
rect 56980 54460 57596 54516
rect 57652 54460 57662 54516
rect 58034 54460 58044 54516
rect 58100 54460 58492 54516
rect 58548 54460 58558 54516
rect 62132 54460 66892 54516
rect 66948 54460 66958 54516
rect 67116 54460 79436 54516
rect 79492 54460 79502 54516
rect 88498 54460 88508 54516
rect 88564 54460 89628 54516
rect 89684 54460 89694 54516
rect 50204 54404 50260 54460
rect 67116 54404 67172 54460
rect 33506 54348 33516 54404
rect 33572 54348 40348 54404
rect 40404 54348 41804 54404
rect 41860 54348 41870 54404
rect 47058 54348 47068 54404
rect 47124 54348 47964 54404
rect 48020 54348 50260 54404
rect 50866 54348 50876 54404
rect 50932 54348 54348 54404
rect 54404 54348 62748 54404
rect 62804 54348 62814 54404
rect 62962 54348 62972 54404
rect 63028 54348 67172 54404
rect 67442 54348 67452 54404
rect 67508 54348 68124 54404
rect 68180 54348 68190 54404
rect 69122 54348 69132 54404
rect 69188 54348 69692 54404
rect 69748 54348 69758 54404
rect 70140 54348 70476 54404
rect 70532 54348 70542 54404
rect 72594 54348 72604 54404
rect 72660 54348 84812 54404
rect 84868 54348 84878 54404
rect 119200 54376 119800 54572
rect 54572 54292 54628 54348
rect 62972 54292 63028 54348
rect 70140 54292 70196 54348
rect 50194 54236 50204 54292
rect 50260 54236 51212 54292
rect 51268 54236 51278 54292
rect 51426 54236 51436 54292
rect 51492 54236 51772 54292
rect 51828 54236 51838 54292
rect 54562 54236 54572 54292
rect 54628 54236 54638 54292
rect 57810 54236 57820 54292
rect 57876 54236 61740 54292
rect 61796 54236 63028 54292
rect 65090 54236 65100 54292
rect 65156 54236 66388 54292
rect 70130 54236 70140 54292
rect 70196 54236 70206 54292
rect 73892 54236 101612 54292
rect 101668 54236 101678 54292
rect 66332 54180 66388 54236
rect 73892 54180 73948 54236
rect 48402 54124 48412 54180
rect 48468 54124 52108 54180
rect 52164 54124 52174 54180
rect 59042 54124 59052 54180
rect 59108 54124 59836 54180
rect 59892 54124 59902 54180
rect 66332 54124 73948 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 51538 54012 51548 54068
rect 51604 54012 51884 54068
rect 51940 54012 53116 54068
rect 53172 54012 53182 54068
rect 53442 54012 53452 54068
rect 53508 54012 62188 54068
rect 66546 54012 66556 54068
rect 66612 54012 67340 54068
rect 67396 54012 67406 54068
rect 46834 53900 46844 53956
rect 46900 53900 49644 53956
rect 49700 53900 49710 53956
rect 59602 53900 59612 53956
rect 59668 53900 60732 53956
rect 60788 53900 60798 53956
rect 62132 53844 62188 54012
rect 66322 53900 66332 53956
rect 66388 53900 67004 53956
rect 67060 53900 67070 53956
rect 42466 53788 42476 53844
rect 42532 53788 43372 53844
rect 43428 53788 43438 53844
rect 48178 53788 48188 53844
rect 48244 53788 48412 53844
rect 48468 53788 48478 53844
rect 48738 53788 48748 53844
rect 48804 53788 49756 53844
rect 49812 53788 49822 53844
rect 51538 53788 51548 53844
rect 51604 53788 52332 53844
rect 52388 53788 52398 53844
rect 57922 53788 57932 53844
rect 57988 53788 59276 53844
rect 59332 53788 59342 53844
rect 59826 53788 59836 53844
rect 59892 53788 60508 53844
rect 60564 53788 60574 53844
rect 62132 53788 68908 53844
rect 68964 53788 68974 53844
rect 45938 53676 45948 53732
rect 46004 53676 47404 53732
rect 47460 53676 47470 53732
rect 49420 53676 50652 53732
rect 50708 53676 50718 53732
rect 50978 53676 50988 53732
rect 51044 53676 51996 53732
rect 52052 53676 52780 53732
rect 52836 53676 52846 53732
rect 59714 53676 59724 53732
rect 59780 53676 61404 53732
rect 61460 53676 62412 53732
rect 62468 53676 62478 53732
rect 62626 53676 62636 53732
rect 62692 53676 63308 53732
rect 63364 53676 65436 53732
rect 65492 53676 65502 53732
rect 67442 53676 67452 53732
rect 67508 53676 70028 53732
rect 70084 53676 71260 53732
rect 71316 53676 71326 53732
rect 31892 53564 45388 53620
rect 45444 53564 49196 53620
rect 49252 53564 49262 53620
rect 31892 53508 31948 53564
rect 49420 53508 49476 53676
rect 30370 53452 30380 53508
rect 30436 53452 31948 53508
rect 47282 53452 47292 53508
rect 47348 53452 48860 53508
rect 48916 53452 49476 53508
rect 50372 53564 50540 53620
rect 50596 53564 50764 53620
rect 50820 53564 51772 53620
rect 51828 53564 51838 53620
rect 57810 53564 57820 53620
rect 57876 53564 58716 53620
rect 58772 53564 62188 53620
rect 62244 53564 65660 53620
rect 65716 53564 65726 53620
rect 50372 53396 50428 53564
rect 50642 53452 50652 53508
rect 50708 53452 51044 53508
rect 51314 53452 51324 53508
rect 51380 53452 52892 53508
rect 52948 53452 52958 53508
rect 55458 53452 55468 53508
rect 55524 53452 56252 53508
rect 56308 53452 56318 53508
rect 58454 53452 58492 53508
rect 58548 53452 58558 53508
rect 62514 53452 62524 53508
rect 62580 53452 63532 53508
rect 63588 53452 66444 53508
rect 66500 53452 66510 53508
rect 68226 53452 68236 53508
rect 68292 53452 70924 53508
rect 70980 53452 104972 53508
rect 105028 53452 105038 53508
rect 47618 53340 47628 53396
rect 47684 53340 49084 53396
rect 49140 53340 50428 53396
rect 50988 53396 51044 53452
rect 50988 53340 51660 53396
rect 51716 53340 51726 53396
rect 53554 53340 53564 53396
rect 53620 53340 62188 53396
rect 62402 53340 62412 53396
rect 62468 53340 66220 53396
rect 66276 53340 77868 53396
rect 77924 53340 77934 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 62132 53284 62188 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 111986 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112270 53340
rect 200 53032 800 53256
rect 47170 53228 47180 53284
rect 47236 53228 48076 53284
rect 48132 53228 48142 53284
rect 52658 53228 52668 53284
rect 52724 53228 53452 53284
rect 53508 53228 54684 53284
rect 54740 53228 54750 53284
rect 58146 53228 58156 53284
rect 58212 53228 61852 53284
rect 61908 53228 61918 53284
rect 62132 53228 67004 53284
rect 67060 53228 67070 53284
rect 54002 53116 54012 53172
rect 54068 53116 56924 53172
rect 56980 53116 56990 53172
rect 57698 53116 57708 53172
rect 57764 53116 58380 53172
rect 58436 53116 58446 53172
rect 58818 53116 58828 53172
rect 58884 53116 59388 53172
rect 59444 53116 59454 53172
rect 60508 53116 62076 53172
rect 62132 53116 62142 53172
rect 64194 53116 64204 53172
rect 64260 53116 68012 53172
rect 68068 53116 69244 53172
rect 69300 53116 69310 53172
rect 60508 53060 60564 53116
rect 51874 53004 51884 53060
rect 51940 53004 54348 53060
rect 54404 53004 54796 53060
rect 54852 53004 54862 53060
rect 56812 53004 59500 53060
rect 59556 53004 60508 53060
rect 60564 53004 60574 53060
rect 61404 53004 70588 53060
rect 70644 53004 70654 53060
rect 119200 53032 119800 53256
rect 56812 52948 56868 53004
rect 61404 52948 61460 53004
rect 49970 52892 49980 52948
rect 50036 52892 53676 52948
rect 53732 52892 53742 52948
rect 55234 52892 55244 52948
rect 55300 52892 56812 52948
rect 56868 52892 56878 52948
rect 58706 52892 58716 52948
rect 58772 52892 61404 52948
rect 61460 52892 61470 52948
rect 61628 52892 66332 52948
rect 66388 52892 66398 52948
rect 53190 52780 53228 52836
rect 53284 52780 57372 52836
rect 57428 52780 57438 52836
rect 57698 52780 57708 52836
rect 57764 52780 59276 52836
rect 59332 52780 59342 52836
rect 61628 52724 61684 52892
rect 62066 52780 62076 52836
rect 62132 52780 63308 52836
rect 63364 52780 63756 52836
rect 63812 52780 63822 52836
rect 69682 52780 69692 52836
rect 69748 52780 70700 52836
rect 70756 52780 72156 52836
rect 72212 52780 72222 52836
rect 108210 52780 108220 52836
rect 108276 52780 114940 52836
rect 114996 52780 115006 52836
rect 48066 52668 48076 52724
rect 48132 52668 52220 52724
rect 52276 52668 52286 52724
rect 52770 52668 52780 52724
rect 52836 52668 56700 52724
rect 56756 52668 61684 52724
rect 47730 52556 47740 52612
rect 47796 52556 50428 52612
rect 50484 52556 50494 52612
rect 51762 52556 51772 52612
rect 51828 52556 54012 52612
rect 54068 52556 54078 52612
rect 57922 52556 57932 52612
rect 57988 52556 58604 52612
rect 58660 52556 60060 52612
rect 60116 52556 60126 52612
rect 60284 52556 63084 52612
rect 63140 52556 63150 52612
rect 116274 52556 116284 52612
rect 116340 52556 116844 52612
rect 116900 52584 119336 52612
rect 116900 52556 119800 52584
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 60284 52500 60340 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 47058 52444 47068 52500
rect 47124 52444 48412 52500
rect 48468 52444 48478 52500
rect 48626 52444 48636 52500
rect 48692 52444 51996 52500
rect 52052 52444 52062 52500
rect 52994 52444 53004 52500
rect 53060 52444 58044 52500
rect 58100 52444 58110 52500
rect 58370 52444 58380 52500
rect 58436 52444 60340 52500
rect 61842 52444 61852 52500
rect 61908 52444 62524 52500
rect 62580 52444 62590 52500
rect 47954 52332 47964 52388
rect 48020 52332 49196 52388
rect 49252 52332 49262 52388
rect 52210 52332 52220 52388
rect 52276 52332 53676 52388
rect 53732 52332 53742 52388
rect 54786 52332 54796 52388
rect 54852 52332 55916 52388
rect 55972 52332 55982 52388
rect 57250 52332 57260 52388
rect 57316 52332 58828 52388
rect 58884 52332 58894 52388
rect 60274 52332 60284 52388
rect 60340 52332 60956 52388
rect 61012 52332 61516 52388
rect 61572 52332 61582 52388
rect 62402 52332 62412 52388
rect 62468 52332 63420 52388
rect 63476 52332 63486 52388
rect 64978 52332 64988 52388
rect 65044 52332 65884 52388
rect 65940 52332 65950 52388
rect 66658 52332 66668 52388
rect 66724 52332 69692 52388
rect 69748 52332 69758 52388
rect 119200 52360 119800 52556
rect 46050 52220 46060 52276
rect 46116 52220 47852 52276
rect 47908 52220 47918 52276
rect 48402 52220 48412 52276
rect 48468 52220 57316 52276
rect 64418 52220 64428 52276
rect 64484 52220 67452 52276
rect 67508 52220 68460 52276
rect 68516 52220 68526 52276
rect 70242 52220 70252 52276
rect 70308 52220 70700 52276
rect 70756 52220 73276 52276
rect 73332 52220 74060 52276
rect 74116 52220 74126 52276
rect 31042 52108 31052 52164
rect 31108 52108 33516 52164
rect 33572 52108 33582 52164
rect 47702 52108 47740 52164
rect 47796 52108 47806 52164
rect 48066 52108 48076 52164
rect 48132 52108 48636 52164
rect 48692 52108 48702 52164
rect 49634 52108 49644 52164
rect 49700 52108 54460 52164
rect 54516 52108 54526 52164
rect 57260 52052 57316 52220
rect 64530 52108 64540 52164
rect 64596 52108 64606 52164
rect 67666 52108 67676 52164
rect 67732 52108 69244 52164
rect 69300 52108 69310 52164
rect 64540 52052 64596 52108
rect 3378 51996 3388 52052
rect 3444 51996 42028 52052
rect 42084 51996 43148 52052
rect 43204 51996 43214 52052
rect 43362 51996 43372 52052
rect 43428 51996 56252 52052
rect 56308 51996 57036 52052
rect 57092 51996 57102 52052
rect 57260 51996 59388 52052
rect 59444 51996 62300 52052
rect 62356 51996 62366 52052
rect 64540 51996 64988 52052
rect 65044 51996 65054 52052
rect 65426 51996 65436 52052
rect 65492 51996 66780 52052
rect 66836 51996 100044 52052
rect 100100 51996 100110 52052
rect 200 51716 800 51912
rect 49942 51884 49980 51940
rect 50036 51884 50046 51940
rect 50306 51884 50316 51940
rect 50372 51884 50988 51940
rect 51044 51884 51054 51940
rect 55682 51884 55692 51940
rect 55748 51884 56364 51940
rect 56420 51884 58828 51940
rect 58884 51884 58894 51940
rect 59154 51884 59164 51940
rect 59220 51884 62188 51940
rect 62244 51884 63084 51940
rect 63140 51884 63150 51940
rect 53890 51772 53900 51828
rect 53956 51772 54908 51828
rect 54964 51772 56476 51828
rect 56532 51772 56542 51828
rect 58930 51772 58940 51828
rect 58996 51772 60396 51828
rect 60452 51772 60462 51828
rect 67218 51772 67228 51828
rect 67284 51772 68572 51828
rect 68628 51772 68638 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 111986 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112270 51772
rect 200 51688 1820 51716
rect 728 51660 1820 51688
rect 1876 51660 1886 51716
rect 50988 51660 51100 51716
rect 51156 51660 51436 51716
rect 51492 51660 55468 51716
rect 55524 51660 55534 51716
rect 64866 51660 64876 51716
rect 64932 51660 65212 51716
rect 65268 51660 66220 51716
rect 66276 51660 72100 51716
rect 50988 51604 51044 51660
rect 72044 51604 72100 51660
rect 29362 51548 29372 51604
rect 29428 51548 49644 51604
rect 49700 51548 49710 51604
rect 50418 51548 50428 51604
rect 50484 51548 51044 51604
rect 51650 51548 51660 51604
rect 51716 51548 53340 51604
rect 53396 51548 53900 51604
rect 53956 51548 59724 51604
rect 59780 51548 59790 51604
rect 66546 51548 66556 51604
rect 66612 51548 67004 51604
rect 67060 51548 67564 51604
rect 67620 51548 68572 51604
rect 68628 51548 68638 51604
rect 72034 51548 72044 51604
rect 72100 51548 73276 51604
rect 73332 51548 73342 51604
rect 31892 51436 45052 51492
rect 45108 51436 45388 51492
rect 45444 51436 47516 51492
rect 47572 51436 47582 51492
rect 49074 51436 49084 51492
rect 49140 51436 50876 51492
rect 50932 51436 51436 51492
rect 51492 51436 51502 51492
rect 55346 51436 55356 51492
rect 55412 51436 56140 51492
rect 56196 51436 56700 51492
rect 56756 51436 57484 51492
rect 57540 51436 57550 51492
rect 57698 51436 57708 51492
rect 57764 51436 58604 51492
rect 58660 51436 58670 51492
rect 68002 51436 68012 51492
rect 68068 51436 69468 51492
rect 69524 51436 78988 51492
rect 31892 51268 31948 51436
rect 78932 51380 78988 51436
rect 45826 51324 45836 51380
rect 45892 51324 46396 51380
rect 46452 51324 46462 51380
rect 48738 51324 48748 51380
rect 48804 51324 59948 51380
rect 60004 51324 60284 51380
rect 60340 51324 60620 51380
rect 60676 51324 62636 51380
rect 62692 51324 63868 51380
rect 63924 51324 65212 51380
rect 65268 51324 65278 51380
rect 65874 51324 65884 51380
rect 65940 51324 68124 51380
rect 68180 51324 68190 51380
rect 68898 51324 68908 51380
rect 68964 51324 69916 51380
rect 69972 51324 69982 51380
rect 71474 51324 71484 51380
rect 71540 51324 72156 51380
rect 72212 51324 72222 51380
rect 72370 51324 72380 51380
rect 72436 51324 73500 51380
rect 73556 51324 73566 51380
rect 78932 51324 91532 51380
rect 91588 51324 91598 51380
rect 17602 51212 17612 51268
rect 17668 51212 31948 51268
rect 45500 51212 48076 51268
rect 48132 51212 48300 51268
rect 48356 51212 48366 51268
rect 49746 51212 49756 51268
rect 49812 51212 50428 51268
rect 50484 51212 50494 51268
rect 53890 51212 53900 51268
rect 53956 51212 54908 51268
rect 54964 51212 54974 51268
rect 56914 51212 56924 51268
rect 56980 51212 70476 51268
rect 70532 51212 71148 51268
rect 71204 51212 71214 51268
rect 45500 51156 45556 51212
rect 34402 51100 34412 51156
rect 34468 51100 34636 51156
rect 34692 51100 45500 51156
rect 45556 51100 45566 51156
rect 46946 51100 46956 51156
rect 47012 51100 50540 51156
rect 50596 51100 52444 51156
rect 52500 51100 52510 51156
rect 63970 51100 63980 51156
rect 64036 51100 65100 51156
rect 65156 51100 65166 51156
rect 73714 51100 73724 51156
rect 73780 51100 100268 51156
rect 100324 51100 100334 51156
rect 48962 50988 48972 51044
rect 49028 50988 50876 51044
rect 50932 50988 52220 51044
rect 52276 50988 53564 51044
rect 53620 50988 53630 51044
rect 55458 50988 55468 51044
rect 55524 50988 62188 51044
rect 64530 50988 64540 51044
rect 64596 50988 64876 51044
rect 64932 50988 64942 51044
rect 119200 51016 119800 51240
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 62132 50932 62188 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 46050 50876 46060 50932
rect 46116 50876 49084 50932
rect 49140 50876 49150 50932
rect 53778 50876 53788 50932
rect 53844 50876 55916 50932
rect 55972 50876 56476 50932
rect 56532 50876 59164 50932
rect 59220 50876 59230 50932
rect 62132 50876 65828 50932
rect 65772 50820 65828 50876
rect 54786 50764 54796 50820
rect 54852 50764 55356 50820
rect 55412 50764 57708 50820
rect 57764 50764 58492 50820
rect 58548 50764 61852 50820
rect 61908 50764 61918 50820
rect 62066 50764 62076 50820
rect 62132 50764 63980 50820
rect 64036 50764 64046 50820
rect 65062 50764 65100 50820
rect 65156 50764 65166 50820
rect 65772 50764 67116 50820
rect 67172 50764 68684 50820
rect 68740 50764 68750 50820
rect 52658 50652 52668 50708
rect 52724 50652 53900 50708
rect 53956 50652 53966 50708
rect 54226 50652 54236 50708
rect 54292 50652 54908 50708
rect 54964 50652 54974 50708
rect 58818 50652 58828 50708
rect 58884 50652 59388 50708
rect 59444 50652 59454 50708
rect 61618 50652 61628 50708
rect 61684 50652 63196 50708
rect 63252 50652 63262 50708
rect 63746 50652 63756 50708
rect 63812 50652 65436 50708
rect 65492 50652 67228 50708
rect 67284 50652 76972 50708
rect 77028 50652 77038 50708
rect 200 50344 800 50568
rect 45826 50540 45836 50596
rect 45892 50540 48300 50596
rect 48356 50540 48748 50596
rect 48804 50540 48814 50596
rect 49410 50540 49420 50596
rect 49476 50540 50428 50596
rect 50866 50540 50876 50596
rect 50932 50540 50942 50596
rect 51174 50540 51212 50596
rect 51268 50540 51278 50596
rect 53778 50540 53788 50596
rect 53844 50540 54572 50596
rect 54628 50540 54638 50596
rect 59938 50540 59948 50596
rect 60004 50540 62188 50596
rect 62244 50540 62254 50596
rect 64316 50540 64988 50596
rect 65044 50540 65660 50596
rect 65716 50540 65726 50596
rect 67778 50540 67788 50596
rect 67844 50540 73948 50596
rect 50372 50484 50428 50540
rect 50876 50484 50932 50540
rect 64316 50484 64372 50540
rect 67788 50484 67844 50540
rect 73892 50484 73948 50540
rect 46386 50428 46396 50484
rect 46452 50428 50204 50484
rect 50260 50428 50270 50484
rect 50372 50428 51940 50484
rect 59490 50428 59500 50484
rect 59556 50428 61628 50484
rect 61684 50428 61694 50484
rect 61842 50428 61852 50484
rect 61908 50428 64316 50484
rect 64372 50428 64382 50484
rect 64764 50428 67844 50484
rect 69906 50428 69916 50484
rect 69972 50428 72268 50484
rect 72324 50428 72334 50484
rect 73892 50428 90188 50484
rect 90244 50428 90254 50484
rect 51884 50372 51940 50428
rect 64764 50372 64820 50428
rect 39554 50316 39564 50372
rect 39620 50316 46396 50372
rect 46452 50316 46462 50372
rect 47954 50316 47964 50372
rect 48020 50316 51660 50372
rect 51716 50316 51726 50372
rect 51884 50316 56812 50372
rect 56868 50316 56878 50372
rect 58370 50316 58380 50372
rect 58436 50316 58828 50372
rect 58884 50316 58894 50372
rect 64754 50316 64764 50372
rect 64820 50316 64830 50372
rect 65314 50316 65324 50372
rect 65380 50316 67676 50372
rect 67732 50316 67742 50372
rect 71698 50316 71708 50372
rect 71764 50316 72716 50372
rect 72772 50316 72782 50372
rect 46834 50204 46844 50260
rect 46900 50204 49308 50260
rect 49364 50204 49374 50260
rect 51762 50204 51772 50260
rect 51828 50204 52332 50260
rect 52388 50204 59500 50260
rect 59556 50204 59566 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 47058 50092 47068 50148
rect 47124 50092 47404 50148
rect 47460 50092 47470 50148
rect 50978 50092 50988 50148
rect 51044 50092 51548 50148
rect 51604 50092 51614 50148
rect 51772 50036 51828 50204
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 111986 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112270 50204
rect 54450 50092 54460 50148
rect 54516 50092 55020 50148
rect 55076 50092 55086 50148
rect 68562 50092 68572 50148
rect 68628 50092 70812 50148
rect 70868 50092 71932 50148
rect 71988 50092 71998 50148
rect 48514 49980 48524 50036
rect 48580 49980 48748 50036
rect 48804 49980 51828 50036
rect 52546 49980 52556 50036
rect 52612 49980 54236 50036
rect 54292 49980 55244 50036
rect 55300 49980 55468 50036
rect 55524 49980 55534 50036
rect 200 49672 800 49896
rect 47394 49868 47404 49924
rect 47460 49868 47852 49924
rect 47908 49868 47918 49924
rect 48850 49868 48860 49924
rect 48916 49868 52108 49924
rect 52164 49868 52174 49924
rect 53666 49868 53676 49924
rect 53732 49868 54012 49924
rect 54068 49868 54348 49924
rect 54404 49868 54414 49924
rect 55122 49868 55132 49924
rect 55188 49868 56364 49924
rect 56420 49868 56430 49924
rect 63410 49868 63420 49924
rect 63476 49868 64204 49924
rect 64260 49868 64270 49924
rect 72258 49868 72268 49924
rect 72324 49868 72492 49924
rect 72548 49868 73164 49924
rect 73220 49868 73230 49924
rect 115490 49868 115500 49924
rect 115556 49896 119336 49924
rect 115556 49868 119800 49896
rect 45490 49756 45500 49812
rect 45556 49756 47068 49812
rect 47124 49756 47134 49812
rect 49746 49756 49756 49812
rect 49812 49756 49980 49812
rect 50036 49756 50046 49812
rect 50372 49756 51884 49812
rect 51940 49756 66276 49812
rect 66434 49756 66444 49812
rect 66500 49756 68124 49812
rect 68180 49756 68190 49812
rect 69794 49756 69804 49812
rect 69860 49756 71484 49812
rect 71540 49756 71550 49812
rect 50372 49700 50428 49756
rect 66220 49700 66276 49756
rect 45266 49644 45276 49700
rect 45332 49644 46732 49700
rect 46788 49644 46798 49700
rect 48402 49644 48412 49700
rect 48468 49644 49196 49700
rect 49252 49644 50428 49700
rect 51538 49644 51548 49700
rect 51604 49644 52556 49700
rect 52612 49644 52622 49700
rect 52770 49644 52780 49700
rect 52836 49644 56252 49700
rect 56308 49644 56318 49700
rect 59042 49644 59052 49700
rect 59108 49644 61292 49700
rect 61348 49644 61358 49700
rect 62850 49644 62860 49700
rect 62916 49644 65324 49700
rect 65380 49644 65390 49700
rect 66220 49644 66780 49700
rect 66836 49644 68572 49700
rect 68628 49644 68638 49700
rect 70354 49644 70364 49700
rect 70420 49644 72268 49700
rect 72324 49644 72334 49700
rect 119200 49672 119800 49868
rect 7522 49532 7532 49588
rect 7588 49532 49532 49588
rect 49588 49532 54236 49588
rect 54292 49532 54302 49588
rect 56802 49532 56812 49588
rect 56868 49532 68348 49588
rect 68404 49532 68414 49588
rect 53218 49420 53228 49476
rect 53284 49420 54684 49476
rect 54740 49420 54750 49476
rect 58818 49420 58828 49476
rect 58884 49420 61068 49476
rect 61124 49420 61134 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 49298 49308 49308 49364
rect 49364 49308 51324 49364
rect 51380 49308 51390 49364
rect 52658 49308 52668 49364
rect 52724 49308 53228 49364
rect 53284 49308 53294 49364
rect 60610 49308 60620 49364
rect 60676 49308 61516 49364
rect 61572 49308 61582 49364
rect 51650 49196 51660 49252
rect 51716 49196 52220 49252
rect 52276 49196 60844 49252
rect 60900 49196 60910 49252
rect 65762 49196 65772 49252
rect 65828 49196 66780 49252
rect 66836 49196 66846 49252
rect 46498 49084 46508 49140
rect 46564 49084 47852 49140
rect 47908 49084 49420 49140
rect 49476 49084 49486 49140
rect 50306 49084 50316 49140
rect 50372 49084 52108 49140
rect 52164 49084 52174 49140
rect 52668 49084 54460 49140
rect 54516 49084 60284 49140
rect 60340 49084 61740 49140
rect 61796 49084 61806 49140
rect 62962 49084 62972 49140
rect 63028 49084 63980 49140
rect 64036 49084 64046 49140
rect 45714 48972 45724 49028
rect 45780 48972 49308 49028
rect 49364 48972 49374 49028
rect 49634 48972 49644 49028
rect 49700 48972 50092 49028
rect 50148 48972 50158 49028
rect 52668 48916 52724 49084
rect 54338 48972 54348 49028
rect 54404 48972 55244 49028
rect 55300 48972 56476 49028
rect 56532 48972 57484 49028
rect 57540 48972 58716 49028
rect 58772 48972 58782 49028
rect 60722 48972 60732 49028
rect 60788 48972 61628 49028
rect 61684 48972 63420 49028
rect 63476 48972 63486 49028
rect 67414 48972 67452 49028
rect 67508 48972 67518 49028
rect 27010 48860 27020 48916
rect 27076 48860 46060 48916
rect 46116 48860 50540 48916
rect 50596 48860 50606 48916
rect 52658 48860 52668 48916
rect 52724 48860 52734 48916
rect 58930 48860 58940 48916
rect 58996 48860 60060 48916
rect 60116 48860 61180 48916
rect 61236 48860 61246 48916
rect 62402 48860 62412 48916
rect 62468 48860 63084 48916
rect 63140 48860 67508 48916
rect 67452 48804 67508 48860
rect 39106 48748 39116 48804
rect 39172 48748 45724 48804
rect 45780 48748 45790 48804
rect 47058 48748 47068 48804
rect 47124 48748 51996 48804
rect 52052 48748 52062 48804
rect 56354 48748 56364 48804
rect 56420 48748 56924 48804
rect 56980 48748 57484 48804
rect 57540 48748 58604 48804
rect 58660 48748 59948 48804
rect 60004 48748 60620 48804
rect 60676 48748 60686 48804
rect 60834 48748 60844 48804
rect 60900 48748 66444 48804
rect 66500 48748 66510 48804
rect 67442 48748 67452 48804
rect 67508 48748 67518 48804
rect 67778 48748 67788 48804
rect 67844 48748 68348 48804
rect 68404 48748 68414 48804
rect 71138 48748 71148 48804
rect 71204 48748 71484 48804
rect 71540 48748 73724 48804
rect 73780 48748 73790 48804
rect 76962 48748 76972 48804
rect 77028 48748 116956 48804
rect 117012 48748 117292 48804
rect 117348 48748 117358 48804
rect 47394 48636 47404 48692
rect 47460 48636 50204 48692
rect 50260 48636 50270 48692
rect 52406 48636 52444 48692
rect 52500 48636 52510 48692
rect 63074 48636 63084 48692
rect 63140 48636 65324 48692
rect 65380 48636 66892 48692
rect 66948 48636 69244 48692
rect 69300 48636 69310 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 111986 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112270 48636
rect 728 48552 1820 48580
rect 200 48524 1820 48552
rect 1876 48524 1886 48580
rect 67414 48524 67452 48580
rect 67508 48524 67518 48580
rect 115490 48524 115500 48580
rect 115556 48552 119336 48580
rect 115556 48524 119800 48552
rect 200 48328 800 48524
rect 43474 48412 43484 48468
rect 43540 48412 57148 48468
rect 57204 48412 58156 48468
rect 58212 48412 58222 48468
rect 61516 48412 64204 48468
rect 64260 48412 64540 48468
rect 64596 48412 64606 48468
rect 14242 48300 14252 48356
rect 14308 48300 31948 48356
rect 45714 48300 45724 48356
rect 45780 48300 47964 48356
rect 48020 48300 48030 48356
rect 49858 48300 49868 48356
rect 49924 48300 53004 48356
rect 53060 48300 53070 48356
rect 31892 48244 31948 48300
rect 61516 48244 61572 48412
rect 61730 48300 61740 48356
rect 61796 48300 63084 48356
rect 63140 48300 63150 48356
rect 67106 48300 67116 48356
rect 67172 48300 68460 48356
rect 68516 48300 68526 48356
rect 119200 48328 119800 48524
rect 31892 48188 52780 48244
rect 52836 48188 52846 48244
rect 55234 48188 55244 48244
rect 55300 48188 57260 48244
rect 57316 48188 57596 48244
rect 57652 48188 61516 48244
rect 61572 48188 61582 48244
rect 62514 48188 62524 48244
rect 62580 48188 62860 48244
rect 62916 48188 62926 48244
rect 63298 48188 63308 48244
rect 63364 48188 63980 48244
rect 64036 48188 64046 48244
rect 68786 48188 68796 48244
rect 68852 48188 70140 48244
rect 70196 48188 70206 48244
rect 46274 48076 46284 48132
rect 46340 48076 48188 48132
rect 48244 48076 48636 48132
rect 48692 48076 48702 48132
rect 50194 48076 50204 48132
rect 50260 48076 50764 48132
rect 50820 48076 50830 48132
rect 53218 48076 53228 48132
rect 53284 48076 54012 48132
rect 54068 48076 54236 48132
rect 54292 48076 56140 48132
rect 56196 48076 56206 48132
rect 56802 48076 56812 48132
rect 56868 48076 57036 48132
rect 57092 48076 58380 48132
rect 58436 48076 58446 48132
rect 60386 48076 60396 48132
rect 60452 48076 61404 48132
rect 61460 48076 61470 48132
rect 61842 48076 61852 48132
rect 61908 48076 63420 48132
rect 63476 48076 64316 48132
rect 64372 48076 64382 48132
rect 65538 48076 65548 48132
rect 65604 48076 66668 48132
rect 66724 48076 66734 48132
rect 67890 48076 67900 48132
rect 67956 48076 69692 48132
rect 69748 48076 80556 48132
rect 80612 48076 80622 48132
rect 56140 48020 56196 48076
rect 48066 47964 48076 48020
rect 48132 47964 54796 48020
rect 54852 47964 54862 48020
rect 56140 47964 62188 48020
rect 63074 47964 63084 48020
rect 63140 47964 65772 48020
rect 65828 47964 65838 48020
rect 66098 47964 66108 48020
rect 66164 47964 67004 48020
rect 67060 47964 67676 48020
rect 67732 47964 67742 48020
rect 54796 47908 54852 47964
rect 62132 47908 62188 47964
rect 54796 47852 56140 47908
rect 56196 47852 61292 47908
rect 61348 47852 61852 47908
rect 61908 47852 61918 47908
rect 62132 47852 63028 47908
rect 115490 47852 115500 47908
rect 115556 47880 119336 47908
rect 115556 47852 119800 47880
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 41234 47740 41244 47796
rect 41300 47740 62524 47796
rect 62580 47740 62590 47796
rect 62972 47684 63028 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 16146 47628 16156 47684
rect 16212 47628 50428 47684
rect 54562 47628 54572 47684
rect 54628 47628 56364 47684
rect 56420 47628 56700 47684
rect 56756 47628 56766 47684
rect 58706 47628 58716 47684
rect 58772 47628 59612 47684
rect 59668 47628 59678 47684
rect 59826 47628 59836 47684
rect 59892 47628 60396 47684
rect 60452 47628 60462 47684
rect 62962 47628 62972 47684
rect 63028 47628 64204 47684
rect 64260 47628 66332 47684
rect 66388 47628 66398 47684
rect 119200 47656 119800 47852
rect 50372 47572 50428 47628
rect 32722 47516 32732 47572
rect 32788 47516 45500 47572
rect 45556 47516 45566 47572
rect 46834 47516 46844 47572
rect 46900 47516 47628 47572
rect 47684 47516 47694 47572
rect 50372 47516 63980 47572
rect 64036 47516 64046 47572
rect 66658 47516 66668 47572
rect 66724 47516 68348 47572
rect 68404 47516 68414 47572
rect 73266 47516 73276 47572
rect 73332 47516 91532 47572
rect 91588 47516 91598 47572
rect 55878 47404 55916 47460
rect 55972 47404 55982 47460
rect 57362 47404 57372 47460
rect 57428 47404 59052 47460
rect 59108 47404 86492 47460
rect 86548 47404 86558 47460
rect 57698 47292 57708 47348
rect 57764 47292 58268 47348
rect 58324 47292 58828 47348
rect 58884 47292 58894 47348
rect 64082 47292 64092 47348
rect 64148 47292 66220 47348
rect 66276 47292 66286 47348
rect 66434 47292 66444 47348
rect 66500 47292 67564 47348
rect 67620 47292 69244 47348
rect 69300 47292 69310 47348
rect 200 46984 800 47208
rect 67778 47180 67788 47236
rect 67844 47180 69804 47236
rect 69860 47180 108332 47236
rect 108388 47180 108398 47236
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 111986 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112270 47068
rect 48962 46956 48972 47012
rect 49028 46956 49532 47012
rect 49588 46956 49598 47012
rect 57586 46956 57596 47012
rect 57652 46956 58716 47012
rect 58772 46956 58782 47012
rect 64306 46956 64316 47012
rect 64372 46956 66668 47012
rect 66724 46956 66734 47012
rect 46834 46844 46844 46900
rect 46900 46844 47292 46900
rect 47348 46844 47358 46900
rect 49858 46844 49868 46900
rect 49924 46844 50428 46900
rect 50484 46844 50494 46900
rect 62290 46844 62300 46900
rect 62356 46844 65772 46900
rect 65828 46844 73276 46900
rect 73332 46844 73342 46900
rect 8418 46732 8428 46788
rect 8484 46732 60844 46788
rect 60900 46732 60910 46788
rect 62132 46732 63196 46788
rect 63252 46732 63532 46788
rect 63588 46732 66220 46788
rect 66276 46732 66286 46788
rect 62132 46676 62188 46732
rect 47618 46620 47628 46676
rect 47684 46620 49868 46676
rect 49924 46620 49934 46676
rect 58146 46620 58156 46676
rect 58212 46620 62188 46676
rect 62962 46620 62972 46676
rect 63028 46620 63756 46676
rect 63812 46620 63822 46676
rect 68002 46620 68012 46676
rect 68068 46620 69020 46676
rect 69076 46620 70364 46676
rect 70420 46620 70430 46676
rect 728 46536 1932 46564
rect 200 46508 1932 46536
rect 1988 46508 1998 46564
rect 53666 46508 53676 46564
rect 53732 46508 54684 46564
rect 54740 46508 55020 46564
rect 55076 46508 57484 46564
rect 57540 46508 57550 46564
rect 58594 46508 58604 46564
rect 58660 46508 59276 46564
rect 59332 46508 59342 46564
rect 63074 46508 63084 46564
rect 63140 46508 67228 46564
rect 67284 46508 108220 46564
rect 108276 46508 108286 46564
rect 118066 46508 118076 46564
rect 118132 46536 119336 46564
rect 118132 46508 119800 46536
rect 200 46312 800 46508
rect 55122 46396 55132 46452
rect 55188 46396 55916 46452
rect 55972 46396 56588 46452
rect 56644 46396 56654 46452
rect 69346 46396 69356 46452
rect 69412 46396 78988 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 78932 46228 78988 46396
rect 119200 46312 119800 46508
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 42914 46172 42924 46228
rect 42980 46172 47740 46228
rect 47796 46172 53452 46228
rect 53508 46172 60844 46228
rect 60900 46172 62188 46228
rect 78932 46172 94892 46228
rect 94948 46172 94958 46228
rect 62132 46116 62188 46172
rect 50306 46060 50316 46116
rect 50372 46060 50652 46116
rect 50708 46060 50718 46116
rect 62132 46060 67452 46116
rect 67508 46060 67518 46116
rect 52210 45948 52220 46004
rect 52276 45948 53900 46004
rect 53956 45948 53966 46004
rect 55346 45948 55356 46004
rect 55412 45948 55692 46004
rect 55748 45948 55758 46004
rect 54114 45836 54124 45892
rect 54180 45836 57932 45892
rect 57988 45836 58604 45892
rect 58660 45836 58670 45892
rect 58930 45836 58940 45892
rect 58996 45836 64092 45892
rect 64148 45836 64158 45892
rect 50866 45724 50876 45780
rect 50932 45724 51436 45780
rect 51492 45724 51502 45780
rect 62850 45724 62860 45780
rect 62916 45724 63868 45780
rect 63924 45724 68012 45780
rect 68068 45724 68078 45780
rect 3042 45612 3052 45668
rect 3108 45612 3500 45668
rect 3556 45612 13412 45668
rect 48402 45612 48412 45668
rect 48468 45612 48972 45668
rect 49028 45612 49196 45668
rect 49252 45612 49980 45668
rect 50036 45612 50204 45668
rect 50260 45612 50270 45668
rect 50372 45612 52220 45668
rect 52276 45612 52286 45668
rect 55346 45612 55356 45668
rect 55412 45612 57260 45668
rect 57316 45612 57596 45668
rect 57652 45612 57662 45668
rect 66994 45612 67004 45668
rect 67060 45612 67564 45668
rect 67620 45612 67630 45668
rect 13356 45332 13412 45612
rect 50372 45556 50428 45612
rect 43586 45500 43596 45556
rect 43652 45500 50428 45556
rect 51202 45500 51212 45556
rect 51268 45500 51548 45556
rect 51604 45500 71372 45556
rect 71428 45500 71438 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 59266 45388 59276 45444
rect 59332 45388 60284 45444
rect 60340 45388 62860 45444
rect 62916 45388 62926 45444
rect 13356 45276 20188 45332
rect 48626 45276 48636 45332
rect 48692 45276 49420 45332
rect 49476 45276 50428 45332
rect 50484 45276 50988 45332
rect 51044 45276 51436 45332
rect 51492 45276 51772 45332
rect 51828 45276 54012 45332
rect 54068 45276 54572 45332
rect 54628 45276 54638 45332
rect 56354 45276 56364 45332
rect 56420 45276 57148 45332
rect 57204 45276 57214 45332
rect 57810 45276 57820 45332
rect 57876 45276 61404 45332
rect 61460 45276 61470 45332
rect 63522 45276 63532 45332
rect 63588 45276 64540 45332
rect 64596 45276 64606 45332
rect 115378 45276 115388 45332
rect 115444 45276 116508 45332
rect 116564 45276 117404 45332
rect 117460 45276 117470 45332
rect 20132 45220 20188 45276
rect 728 45192 1932 45220
rect 200 45164 1932 45192
rect 1988 45164 1998 45220
rect 20132 45164 42140 45220
rect 42196 45164 42206 45220
rect 51986 45164 51996 45220
rect 52052 45164 53228 45220
rect 53284 45164 53676 45220
rect 53732 45164 53742 45220
rect 55794 45164 55804 45220
rect 55860 45164 58828 45220
rect 58884 45164 59388 45220
rect 59444 45164 59454 45220
rect 64204 45164 64316 45220
rect 64372 45164 65772 45220
rect 65828 45164 65838 45220
rect 115490 45164 115500 45220
rect 115556 45192 119336 45220
rect 115556 45164 119800 45192
rect 200 44968 800 45164
rect 41906 45052 41916 45108
rect 41972 45052 45612 45108
rect 45668 45052 46956 45108
rect 47012 45052 47516 45108
rect 47572 45052 47582 45108
rect 57138 45052 57148 45108
rect 57204 45052 58492 45108
rect 58548 45052 58558 45108
rect 58930 45052 58940 45108
rect 58996 45052 59612 45108
rect 59668 45052 61292 45108
rect 61348 45052 61358 45108
rect 64204 44996 64260 45164
rect 53218 44940 53228 44996
rect 53284 44940 53788 44996
rect 53844 44940 55468 44996
rect 55524 44940 55534 44996
rect 55906 44940 55916 44996
rect 55972 44940 58716 44996
rect 58772 44940 58782 44996
rect 61730 44940 61740 44996
rect 61796 44940 64260 44996
rect 65436 45052 68796 45108
rect 68852 45052 68862 45108
rect 65436 44884 65492 45052
rect 119200 44968 119800 45164
rect 29362 44828 29372 44884
rect 29428 44828 38668 44884
rect 54562 44828 54572 44884
rect 54628 44828 55356 44884
rect 55412 44828 55422 44884
rect 58482 44828 58492 44884
rect 58548 44828 59500 44884
rect 59556 44828 60060 44884
rect 60116 44828 60126 44884
rect 62132 44828 65492 44884
rect 65772 44828 66444 44884
rect 66500 44828 67228 44884
rect 67284 44828 67294 44884
rect 80546 44828 80556 44884
rect 80612 44828 115164 44884
rect 115220 44828 115230 44884
rect 38612 44772 38668 44828
rect 62132 44772 62188 44828
rect 38612 44716 54460 44772
rect 54516 44716 55244 44772
rect 55300 44716 55310 44772
rect 55682 44716 55692 44772
rect 55748 44716 62188 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 55692 44660 55748 44716
rect 65772 44660 65828 44828
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 50530 44604 50540 44660
rect 50596 44604 50876 44660
rect 50932 44604 55748 44660
rect 61058 44604 61068 44660
rect 61124 44604 65828 44660
rect 66322 44604 66332 44660
rect 66388 44604 73948 44660
rect 61068 44548 61124 44604
rect 73892 44548 73948 44604
rect 51538 44492 51548 44548
rect 51604 44492 61124 44548
rect 61954 44492 61964 44548
rect 62020 44492 62748 44548
rect 62804 44492 62814 44548
rect 63298 44492 63308 44548
rect 63364 44492 65324 44548
rect 65380 44492 66668 44548
rect 66724 44492 66734 44548
rect 73892 44492 115388 44548
rect 115444 44492 115454 44548
rect 50418 44380 50428 44436
rect 50484 44380 51996 44436
rect 52052 44380 52062 44436
rect 58370 44380 58380 44436
rect 58436 44380 59500 44436
rect 59556 44380 59566 44436
rect 61618 44380 61628 44436
rect 61684 44380 79772 44436
rect 79828 44380 79838 44436
rect 49970 44268 49980 44324
rect 50036 44268 50932 44324
rect 50876 44100 50932 44268
rect 61292 44268 62188 44324
rect 62244 44268 62412 44324
rect 62468 44268 62478 44324
rect 65650 44268 65660 44324
rect 65716 44268 66108 44324
rect 66164 44268 66174 44324
rect 66882 44268 66892 44324
rect 66948 44268 67900 44324
rect 67956 44268 67966 44324
rect 51314 44156 51324 44212
rect 51380 44156 51772 44212
rect 51828 44156 53116 44212
rect 53172 44156 53900 44212
rect 53956 44156 54460 44212
rect 54516 44156 54526 44212
rect 61292 44100 61348 44268
rect 66892 44212 66948 44268
rect 61506 44156 61516 44212
rect 61572 44156 62972 44212
rect 63028 44156 63038 44212
rect 63410 44156 63420 44212
rect 63476 44156 63980 44212
rect 64036 44156 64204 44212
rect 64260 44156 64270 44212
rect 64428 44156 66948 44212
rect 64428 44100 64484 44156
rect 47058 44044 47068 44100
rect 47124 44044 47852 44100
rect 47908 44044 48076 44100
rect 48132 44044 48142 44100
rect 50866 44044 50876 44100
rect 50932 44044 51884 44100
rect 51940 44044 51950 44100
rect 52434 44044 52444 44100
rect 52500 44044 53452 44100
rect 53508 44044 53518 44100
rect 54114 44044 54124 44100
rect 54180 44044 54796 44100
rect 54852 44044 54862 44100
rect 60050 44044 60060 44100
rect 60116 44044 61628 44100
rect 61684 44044 61694 44100
rect 62178 44044 62188 44100
rect 62244 44044 63196 44100
rect 63252 44044 64484 44100
rect 66994 44044 67004 44100
rect 67060 44044 68460 44100
rect 68516 44044 68526 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 200 43624 800 43848
rect 54796 43764 54852 44044
rect 55346 43932 55356 43988
rect 55412 43932 55804 43988
rect 55860 43932 67116 43988
rect 67172 43932 67182 43988
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 55234 43820 55244 43876
rect 55300 43820 57820 43876
rect 57876 43820 57886 43876
rect 61954 43820 61964 43876
rect 62020 43820 63868 43876
rect 63924 43820 63934 43876
rect 64194 43820 64204 43876
rect 64260 43820 64540 43876
rect 64596 43820 66332 43876
rect 66388 43820 66398 43876
rect 53676 43708 53788 43764
rect 53844 43708 53854 43764
rect 54796 43708 55356 43764
rect 55412 43708 57540 43764
rect 60274 43708 60284 43764
rect 60340 43708 62076 43764
rect 62132 43708 62142 43764
rect 62290 43708 62300 43764
rect 62356 43708 63532 43764
rect 63588 43708 63598 43764
rect 63868 43708 65660 43764
rect 65716 43708 65726 43764
rect 67442 43708 67452 43764
rect 67508 43708 68236 43764
rect 68292 43708 118188 43764
rect 118244 43708 118254 43764
rect 53676 43652 53732 43708
rect 57484 43652 57540 43708
rect 63868 43652 63924 43708
rect 49522 43596 49532 43652
rect 49588 43596 50764 43652
rect 50820 43596 52892 43652
rect 52948 43596 53732 43652
rect 54226 43596 54236 43652
rect 54292 43596 55132 43652
rect 55188 43596 55198 43652
rect 57474 43596 57484 43652
rect 57540 43596 59388 43652
rect 59444 43596 61740 43652
rect 61796 43596 61806 43652
rect 63074 43596 63084 43652
rect 63140 43596 63924 43652
rect 119200 43624 119800 43848
rect 59602 43484 59612 43540
rect 59668 43484 60508 43540
rect 60564 43484 60574 43540
rect 61170 43484 61180 43540
rect 61236 43484 62748 43540
rect 62804 43484 65324 43540
rect 65380 43484 65390 43540
rect 10882 43372 10892 43428
rect 10948 43372 48300 43428
rect 48356 43372 49532 43428
rect 49588 43372 49598 43428
rect 54898 43372 54908 43428
rect 54964 43372 56364 43428
rect 56420 43372 56430 43428
rect 61842 43372 61852 43428
rect 61908 43372 63084 43428
rect 63140 43372 63150 43428
rect 73938 43372 73948 43428
rect 74004 43372 75068 43428
rect 75124 43372 82348 43428
rect 82404 43372 82414 43428
rect 87266 43372 87276 43428
rect 87332 43372 87836 43428
rect 87892 43372 100828 43428
rect 100884 43372 100894 43428
rect 101826 43372 101836 43428
rect 101892 43372 114940 43428
rect 114996 43372 115006 43428
rect 59154 43260 59164 43316
rect 59220 43260 59948 43316
rect 60004 43260 60014 43316
rect 62402 43260 62412 43316
rect 62468 43260 64428 43316
rect 64484 43260 65212 43316
rect 65268 43260 65278 43316
rect 41122 43148 41132 43204
rect 41188 43148 53452 43204
rect 53508 43148 53518 43204
rect 116274 43148 116284 43204
rect 116340 43148 116844 43204
rect 116900 43176 119336 43204
rect 116900 43148 119800 43176
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 48850 43036 48860 43092
rect 48916 43036 50428 43092
rect 50484 43036 60060 43092
rect 60116 43036 60620 43092
rect 60676 43036 61292 43092
rect 61348 43036 61358 43092
rect 52210 42924 52220 42980
rect 52276 42924 60508 42980
rect 60564 42924 61516 42980
rect 61572 42924 62188 42980
rect 119200 42952 119800 43148
rect 62132 42868 62188 42924
rect 10546 42812 10556 42868
rect 10612 42812 41916 42868
rect 41972 42812 41982 42868
rect 53442 42812 53452 42868
rect 53508 42812 54908 42868
rect 54964 42812 54974 42868
rect 56354 42812 56364 42868
rect 56420 42812 57932 42868
rect 57988 42812 58716 42868
rect 58772 42812 59948 42868
rect 60004 42812 60014 42868
rect 62132 42812 63980 42868
rect 64036 42812 64046 42868
rect 66770 42812 66780 42868
rect 66836 42812 73948 42868
rect 74004 42812 74014 42868
rect 48178 42700 48188 42756
rect 48244 42700 49868 42756
rect 49924 42700 51772 42756
rect 51828 42700 51838 42756
rect 49746 42588 49756 42644
rect 49812 42588 51548 42644
rect 51604 42588 51614 42644
rect 53666 42588 53676 42644
rect 53732 42588 55692 42644
rect 55748 42588 55758 42644
rect 59378 42588 59388 42644
rect 59444 42588 61404 42644
rect 61460 42588 61470 42644
rect 61618 42588 61628 42644
rect 61684 42588 63532 42644
rect 63588 42588 63598 42644
rect 200 42280 800 42504
rect 15922 42476 15932 42532
rect 15988 42476 47740 42532
rect 47796 42476 51436 42532
rect 51492 42476 51502 42532
rect 56802 42476 56812 42532
rect 56868 42476 58156 42532
rect 58212 42476 59612 42532
rect 59668 42476 59678 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 58146 42028 58156 42084
rect 58212 42028 59164 42084
rect 59220 42028 59230 42084
rect 59378 42028 59388 42084
rect 59444 42028 60172 42084
rect 60228 42028 61852 42084
rect 61908 42028 63980 42084
rect 64036 42028 64046 42084
rect 48300 41916 50876 41972
rect 50932 41916 50942 41972
rect 51874 41916 51884 41972
rect 51940 41916 56364 41972
rect 56420 41916 56430 41972
rect 59826 41916 59836 41972
rect 59892 41916 61180 41972
rect 61236 41916 61246 41972
rect 91522 41916 91532 41972
rect 91588 41916 114380 41972
rect 114436 41916 114940 41972
rect 114996 41916 115006 41972
rect 48300 41860 48356 41916
rect 200 41608 800 41832
rect 44930 41804 44940 41860
rect 44996 41804 48300 41860
rect 48356 41804 48366 41860
rect 49858 41804 49868 41860
rect 49924 41804 52780 41860
rect 52836 41804 53452 41860
rect 53508 41804 53900 41860
rect 53956 41804 54460 41860
rect 54516 41804 54526 41860
rect 115826 41804 115836 41860
rect 115892 41832 119336 41860
rect 115892 41804 119800 41832
rect 37538 41692 37548 41748
rect 37604 41692 48748 41748
rect 48804 41692 52556 41748
rect 52612 41692 52622 41748
rect 119200 41608 119800 41804
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 3266 41244 3276 41300
rect 3332 41244 22652 41300
rect 22708 41244 22718 41300
rect 53554 41244 53564 41300
rect 53620 41244 54236 41300
rect 54292 41244 54302 41300
rect 58258 41244 58268 41300
rect 58324 41244 59500 41300
rect 59556 41244 60284 41300
rect 60340 41244 61180 41300
rect 61236 41244 61404 41300
rect 61460 41244 61470 41300
rect 3602 41132 3612 41188
rect 3668 41132 32732 41188
rect 32788 41132 32798 41188
rect 49410 41132 49420 41188
rect 49476 41132 49868 41188
rect 49924 41132 49934 41188
rect 50372 41132 57372 41188
rect 57428 41132 58492 41188
rect 58548 41132 59052 41188
rect 59108 41132 59118 41188
rect 100818 41132 100828 41188
rect 100884 41132 115276 41188
rect 115332 41132 115342 41188
rect 50372 41076 50428 41132
rect 47628 41020 50428 41076
rect 50530 41020 50540 41076
rect 50596 41020 50988 41076
rect 51044 41020 51054 41076
rect 52658 41020 52668 41076
rect 52724 41020 53564 41076
rect 53620 41020 53630 41076
rect 47628 40964 47684 41020
rect 52668 40964 52724 41020
rect 47618 40908 47628 40964
rect 47684 40908 47694 40964
rect 49186 40908 49196 40964
rect 49252 40908 52724 40964
rect 61618 40908 61628 40964
rect 61684 40908 62748 40964
rect 62804 40908 91868 40964
rect 91924 40908 91934 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 56354 40684 56364 40740
rect 56420 40684 57708 40740
rect 57764 40684 57774 40740
rect 43138 40572 43148 40628
rect 43204 40572 58156 40628
rect 58212 40572 58828 40628
rect 58884 40572 58894 40628
rect 61170 40572 61180 40628
rect 61236 40572 61964 40628
rect 62020 40572 62030 40628
rect 728 40488 1708 40516
rect 200 40460 1708 40488
rect 1764 40460 1774 40516
rect 51538 40460 51548 40516
rect 51604 40460 53676 40516
rect 53732 40460 53742 40516
rect 115490 40460 115500 40516
rect 115556 40488 119336 40516
rect 115556 40460 119800 40488
rect 200 40264 800 40460
rect 32162 40348 32172 40404
rect 32228 40348 37772 40404
rect 37828 40348 37838 40404
rect 48738 40348 48748 40404
rect 48804 40348 49420 40404
rect 49476 40348 49486 40404
rect 61506 40348 61516 40404
rect 61572 40348 62412 40404
rect 62468 40348 101836 40404
rect 101892 40348 101902 40404
rect 36082 40236 36092 40292
rect 36148 40236 45836 40292
rect 45892 40236 47404 40292
rect 47460 40236 47470 40292
rect 55570 40236 55580 40292
rect 55636 40236 56476 40292
rect 56532 40236 56542 40292
rect 58594 40236 58604 40292
rect 58660 40236 60508 40292
rect 60564 40236 60574 40292
rect 62132 40236 102508 40292
rect 119200 40264 119800 40460
rect 56476 40180 56532 40236
rect 62132 40180 62188 40236
rect 56476 40124 62188 40180
rect 102452 40180 102508 40236
rect 102452 40124 116060 40180
rect 116116 40124 116126 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 22642 39788 22652 39844
rect 22708 39788 65548 39844
rect 65604 39788 65614 39844
rect 119200 39732 119800 39816
rect 8754 39676 8764 39732
rect 8820 39676 31948 39732
rect 48402 39676 48412 39732
rect 48468 39676 49644 39732
rect 49700 39676 49868 39732
rect 49924 39676 49934 39732
rect 116274 39676 116284 39732
rect 116340 39676 117068 39732
rect 117124 39676 119800 39732
rect 31892 39620 31948 39676
rect 3042 39564 3052 39620
rect 3108 39564 3612 39620
rect 3668 39564 3678 39620
rect 31892 39564 57596 39620
rect 57652 39564 57662 39620
rect 62962 39564 62972 39620
rect 63028 39564 74060 39620
rect 74116 39564 74126 39620
rect 119200 39592 119800 39676
rect 47394 39452 47404 39508
rect 47460 39452 48972 39508
rect 49028 39452 49038 39508
rect 49186 39452 49196 39508
rect 49252 39452 50204 39508
rect 50260 39452 50428 39508
rect 50372 39396 50428 39452
rect 50372 39340 62636 39396
rect 62692 39340 63420 39396
rect 63476 39340 63486 39396
rect 115602 39228 115612 39284
rect 115668 39228 117292 39284
rect 117348 39228 117358 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 728 39144 1932 39172
rect 200 39116 1932 39144
rect 1988 39116 1998 39172
rect 200 38920 800 39116
rect 62850 38892 62860 38948
rect 62916 38892 63868 38948
rect 63924 38892 63934 38948
rect 118066 38668 118076 38724
rect 118132 38668 118142 38724
rect 118076 38500 118132 38668
rect 118076 38472 119336 38500
rect 118076 38444 119800 38472
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 119200 38248 119800 38444
rect 3378 37884 3388 37940
rect 3444 37884 8428 37940
rect 8484 37884 8494 37940
rect 728 37800 1932 37828
rect 200 37772 1932 37800
rect 1988 37772 1998 37828
rect 3042 37772 3052 37828
rect 3108 37772 3500 37828
rect 3556 37772 55132 37828
rect 55188 37772 56028 37828
rect 56084 37772 56364 37828
rect 56420 37772 56430 37828
rect 68450 37772 68460 37828
rect 68516 37772 103292 37828
rect 103348 37772 103358 37828
rect 103506 37772 103516 37828
rect 103572 37772 114828 37828
rect 114884 37772 114894 37828
rect 200 37576 800 37772
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 53554 37436 53564 37492
rect 53620 37436 54236 37492
rect 54292 37436 54302 37492
rect 54562 37212 54572 37268
rect 54628 37212 56476 37268
rect 56532 37212 56542 37268
rect 728 37128 1932 37156
rect 200 37100 1932 37128
rect 1988 37100 1998 37156
rect 54674 37100 54684 37156
rect 54740 37100 55468 37156
rect 55524 37100 55534 37156
rect 200 36904 800 37100
rect 45938 36988 45948 37044
rect 46004 36988 46620 37044
rect 46676 36988 53564 37044
rect 53620 36988 54908 37044
rect 54964 36988 54974 37044
rect 119200 36904 119800 37128
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 3266 36540 3276 36596
rect 3332 36540 37548 36596
rect 37604 36540 37614 36596
rect 116162 36316 116172 36372
rect 116228 36316 117068 36372
rect 117124 36316 117134 36372
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 728 35784 2156 35812
rect 200 35756 2156 35784
rect 2212 35756 2222 35812
rect 117058 35756 117068 35812
rect 117124 35784 119336 35812
rect 117124 35756 119800 35784
rect 200 35560 800 35756
rect 95666 35644 95676 35700
rect 95732 35644 114492 35700
rect 114548 35644 114940 35700
rect 114996 35644 115006 35700
rect 119200 35560 119800 35756
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 110226 35196 110236 35252
rect 110292 35196 112812 35252
rect 112868 35196 112878 35252
rect 3378 35084 3388 35140
rect 3444 35084 8764 35140
rect 8820 35084 8830 35140
rect 115826 35084 115836 35140
rect 115892 35112 119336 35140
rect 115892 35084 119800 35112
rect 119200 34888 119800 35084
rect 58594 34636 58604 34692
rect 58660 34636 95676 34692
rect 95732 34636 95742 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 728 34440 1932 34468
rect 200 34412 1932 34440
rect 1988 34412 1998 34468
rect 200 34216 800 34412
rect 46050 34188 46060 34244
rect 46116 34188 47180 34244
rect 47236 34188 47246 34244
rect 3042 33964 3052 34020
rect 3108 33964 3612 34020
rect 3668 33964 45052 34020
rect 45108 33964 45118 34020
rect 110002 33964 110012 34020
rect 110068 33964 114604 34020
rect 114660 33964 115164 34020
rect 115220 33964 115230 34020
rect 116050 33964 116060 34020
rect 116116 33964 117180 34020
rect 117236 33964 118076 34020
rect 118132 33964 118142 34020
rect 728 33768 1932 33796
rect 200 33740 1932 33768
rect 1988 33740 1998 33796
rect 200 33544 800 33740
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 119200 33684 119800 33768
rect 115490 33628 115500 33684
rect 115556 33628 119800 33684
rect 94882 33516 94892 33572
rect 94948 33516 112588 33572
rect 112644 33516 112654 33572
rect 119200 33544 119800 33628
rect 37762 33404 37772 33460
rect 37828 33404 46396 33460
rect 46452 33404 47740 33460
rect 47796 33404 48524 33460
rect 48580 33404 48590 33460
rect 46610 33292 46620 33348
rect 46676 33292 48188 33348
rect 48244 33292 48580 33348
rect 48524 33236 48580 33292
rect 45378 33180 45388 33236
rect 45444 33180 46956 33236
rect 47012 33180 47022 33236
rect 48514 33180 48524 33236
rect 48580 33180 48590 33236
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 60060 32844 60396 32900
rect 60452 32844 60462 32900
rect 60060 32788 60116 32844
rect 60050 32732 60060 32788
rect 60116 32732 60126 32788
rect 102452 32620 114940 32676
rect 114996 32620 116620 32676
rect 116676 32620 116686 32676
rect 102452 32452 102508 32620
rect 200 32228 800 32424
rect 3266 32396 3276 32452
rect 3332 32396 36204 32452
rect 36260 32396 36270 32452
rect 95218 32396 95228 32452
rect 95284 32396 102508 32452
rect 112578 32284 112588 32340
rect 112644 32284 115388 32340
rect 115444 32284 116396 32340
rect 116452 32284 116462 32340
rect 200 32200 1932 32228
rect 728 32172 1932 32200
rect 1988 32172 1998 32228
rect 119200 32200 119800 32424
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 48178 31948 48188 32004
rect 48244 31948 48412 32004
rect 48468 31948 58828 32004
rect 58884 31948 60620 32004
rect 60676 31948 60686 32004
rect 119200 31528 119800 31752
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 12338 31164 12348 31220
rect 12404 31164 34636 31220
rect 34692 31164 34702 31220
rect 200 30856 800 31080
rect 34402 31052 34412 31108
rect 34468 31052 57148 31108
rect 57204 31052 57214 31108
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 115490 30380 115500 30436
rect 115556 30408 119336 30436
rect 115556 30380 119800 30408
rect 3378 30156 3388 30212
rect 3444 30156 15932 30212
rect 15988 30156 15998 30212
rect 114370 30156 114380 30212
rect 114436 30156 115500 30212
rect 115556 30156 115566 30212
rect 119200 30184 119800 30380
rect 67554 30044 67564 30100
rect 67620 30044 72268 30100
rect 72324 30044 76524 30100
rect 76580 30044 76590 30100
rect 69346 29932 69356 29988
rect 69412 29932 75068 29988
rect 75124 29932 75134 29988
rect 114930 29932 114940 29988
rect 114996 29932 116284 29988
rect 116340 29932 117404 29988
rect 117460 29932 117470 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 200 29652 800 29736
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 200 29512 800 29596
rect 200 28840 800 29064
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 119200 28840 119800 29064
rect 68114 28588 68124 28644
rect 68180 28588 70252 28644
rect 70308 28588 70318 28644
rect 47730 28476 47740 28532
rect 47796 28476 48300 28532
rect 48356 28476 49420 28532
rect 49476 28476 49486 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 200 27496 800 27720
rect 71362 27692 71372 27748
rect 71428 27692 84140 27748
rect 84196 27692 84206 27748
rect 119200 27496 119800 27720
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 3378 27244 3388 27300
rect 3444 27244 7532 27300
rect 7588 27244 7598 27300
rect 31892 27244 46060 27300
rect 46116 27244 47292 27300
rect 47348 27244 47358 27300
rect 31892 27076 31948 27244
rect 46834 27132 46844 27188
rect 46900 27132 47852 27188
rect 47908 27132 48300 27188
rect 48356 27132 48366 27188
rect 9650 27020 9660 27076
rect 9716 27020 31948 27076
rect 115490 27020 115500 27076
rect 115556 27048 119336 27076
rect 115556 27020 119800 27048
rect 29474 26908 29484 26964
rect 29540 26908 44716 26964
rect 44772 26908 46620 26964
rect 46676 26908 46686 26964
rect 116162 26908 116172 26964
rect 116228 26908 117068 26964
rect 117124 26908 117134 26964
rect 119200 26824 119800 27020
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 62738 26460 62748 26516
rect 62804 26460 63196 26516
rect 63252 26460 69356 26516
rect 69412 26460 69422 26516
rect 728 26376 1708 26404
rect 200 26348 1708 26376
rect 1764 26348 1774 26404
rect 200 26152 800 26348
rect 80098 26236 80108 26292
rect 80164 26236 114380 26292
rect 114436 26236 114940 26292
rect 114996 26236 115006 26292
rect 70802 26012 70812 26068
rect 70868 26012 72380 26068
rect 72436 26012 72446 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 69458 25788 69468 25844
rect 69524 25788 70924 25844
rect 70980 25788 70990 25844
rect 3378 25676 3388 25732
rect 3444 25676 5852 25732
rect 5908 25676 5918 25732
rect 115826 25676 115836 25732
rect 115892 25704 119336 25732
rect 115892 25676 119800 25704
rect 119200 25480 119800 25676
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 728 25032 1932 25060
rect 200 25004 1932 25032
rect 1988 25004 1998 25060
rect 200 24808 800 25004
rect 79762 24892 79772 24948
rect 79828 24892 86940 24948
rect 86996 24892 87006 24948
rect 3042 24556 3052 24612
rect 3108 24556 3500 24612
rect 3556 24556 17612 24612
rect 17668 24556 17678 24612
rect 86482 24444 86492 24500
rect 86548 24444 114716 24500
rect 114772 24444 114782 24500
rect 728 24360 1932 24388
rect 200 24332 1932 24360
rect 1988 24332 1998 24388
rect 200 24136 800 24332
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 119200 24136 119800 24360
rect 17826 23884 17836 23940
rect 17892 23884 46060 23940
rect 46116 23884 47460 23940
rect 47404 23828 47460 23884
rect 31892 23772 44716 23828
rect 44772 23772 46620 23828
rect 46676 23772 46686 23828
rect 47394 23772 47404 23828
rect 47460 23772 60172 23828
rect 60228 23772 63868 23828
rect 63924 23772 63934 23828
rect 31892 23716 31948 23772
rect 26114 23660 26124 23716
rect 26180 23660 31948 23716
rect 46834 23660 46844 23716
rect 46900 23660 47852 23716
rect 47908 23660 48524 23716
rect 48580 23660 78316 23716
rect 78372 23660 79100 23716
rect 79156 23660 79166 23716
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 77634 23100 77644 23156
rect 77700 23100 78540 23156
rect 78596 23100 78606 23156
rect 728 23016 1932 23044
rect 200 22988 1932 23016
rect 1988 22988 1998 23044
rect 3042 22988 3052 23044
rect 3108 22988 3500 23044
rect 3556 22988 12348 23044
rect 12404 22988 12414 23044
rect 200 22792 800 22988
rect 119200 22792 119800 23016
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 47170 22428 47180 22484
rect 47236 22428 48188 22484
rect 48244 22428 48524 22484
rect 48580 22428 48590 22484
rect 76514 22316 76524 22372
rect 76580 22316 77532 22372
rect 77588 22316 77598 22372
rect 115490 22316 115500 22372
rect 115556 22344 119336 22372
rect 115556 22316 119800 22344
rect 46386 22204 46396 22260
rect 46452 22204 46844 22260
rect 46900 22204 47740 22260
rect 47796 22204 59836 22260
rect 59892 22204 59902 22260
rect 4386 22092 4396 22148
rect 4452 22092 26012 22148
rect 26068 22092 26078 22148
rect 44258 22092 44268 22148
rect 44324 22092 46060 22148
rect 46116 22092 46126 22148
rect 48514 22092 48524 22148
rect 48580 22092 68796 22148
rect 68852 22092 68862 22148
rect 119200 22120 119800 22316
rect 45042 21980 45052 22036
rect 45108 21980 45500 22036
rect 45556 21980 46956 22036
rect 47012 21980 47022 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 200 21476 800 21672
rect 44482 21644 44492 21700
rect 44548 21644 47180 21700
rect 47236 21644 47246 21700
rect 90692 21532 91308 21588
rect 91364 21532 110012 21588
rect 110068 21532 110078 21588
rect 200 21448 1820 21476
rect 728 21420 1820 21448
rect 1876 21420 1886 21476
rect 34514 21420 34524 21476
rect 34580 21420 45052 21476
rect 45108 21420 45118 21476
rect 77522 21420 77532 21476
rect 77588 21420 90636 21476
rect 90692 21420 90748 21532
rect 93090 21420 93100 21476
rect 93156 21420 94108 21476
rect 94164 21420 95004 21476
rect 95060 21420 95070 21476
rect 3042 21308 3052 21364
rect 3108 21308 3612 21364
rect 3668 21308 39452 21364
rect 39508 21308 39518 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 728 21000 1932 21028
rect 200 20972 1932 21000
rect 1988 20972 1998 21028
rect 115154 20972 115164 21028
rect 115220 21000 119336 21028
rect 115220 20972 119800 21000
rect 200 20776 800 20972
rect 39778 20860 39788 20916
rect 39844 20860 40236 20916
rect 40292 20860 41132 20916
rect 41188 20860 41198 20916
rect 45826 20860 45836 20916
rect 45892 20860 47628 20916
rect 47684 20860 47694 20916
rect 48290 20860 48300 20916
rect 48356 20860 48972 20916
rect 49028 20860 49038 20916
rect 90514 20748 90524 20804
rect 90580 20748 91532 20804
rect 91588 20748 91598 20804
rect 92194 20748 92204 20804
rect 92260 20748 95228 20804
rect 95284 20748 95294 20804
rect 119200 20776 119800 20972
rect 92306 20636 92316 20692
rect 92372 20636 93100 20692
rect 93156 20636 93166 20692
rect 68786 20524 68796 20580
rect 68852 20524 90076 20580
rect 90132 20524 92204 20580
rect 92260 20524 92270 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 45490 20076 45500 20132
rect 45556 20076 46620 20132
rect 46676 20076 46956 20132
rect 47012 20076 47022 20132
rect 47170 19964 47180 20020
rect 47236 19964 48300 20020
rect 48356 19964 48366 20020
rect 5618 19740 5628 19796
rect 5684 19740 46396 19796
rect 46452 19740 47516 19796
rect 47572 19740 47740 19796
rect 47796 19740 47806 19796
rect 200 19432 800 19656
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 119200 19432 119800 19656
rect 115490 18956 115500 19012
rect 115556 18984 119336 19012
rect 115556 18956 119800 18984
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 119200 18760 119800 18956
rect 728 18312 1820 18340
rect 200 18284 1820 18312
rect 1876 18284 1886 18340
rect 200 18088 800 18284
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 84802 17612 84812 17668
rect 84868 17612 112364 17668
rect 112420 17612 112430 17668
rect 119200 17416 119800 17640
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 728 16968 1820 16996
rect 200 16940 1820 16968
rect 1876 16940 1886 16996
rect 118066 16940 118076 16996
rect 118132 16940 119364 16996
rect 200 16744 800 16940
rect 3042 16828 3052 16884
rect 3108 16828 3500 16884
rect 3556 16828 13580 16884
rect 13636 16828 13646 16884
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 119308 16436 119364 16940
rect 119084 16380 119364 16436
rect 119084 16324 119140 16380
rect 728 16296 1932 16324
rect 200 16268 1932 16296
rect 1988 16268 1998 16324
rect 119084 16296 119336 16324
rect 119084 16268 119800 16296
rect 200 16072 800 16268
rect 119200 16072 119800 16268
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 54450 15372 54460 15428
rect 54516 15372 114492 15428
rect 114548 15372 114940 15428
rect 114996 15372 115006 15428
rect 13570 15148 13580 15204
rect 13636 15148 53676 15204
rect 53732 15148 54124 15204
rect 54180 15148 54190 15204
rect 200 14728 800 14952
rect 115826 14924 115836 14980
rect 115892 14952 119336 14980
rect 115892 14924 119800 14952
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 119200 14728 119800 14924
rect 102452 14476 114492 14532
rect 114548 14476 114940 14532
rect 114996 14476 115006 14532
rect 102452 14308 102508 14476
rect 100258 14252 100268 14308
rect 100324 14252 102508 14308
rect 115826 14252 115836 14308
rect 115892 14280 119336 14308
rect 115892 14252 119800 14280
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 119200 14056 119800 14252
rect 200 13384 800 13608
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 19618 12684 19628 12740
rect 19684 12684 29372 12740
rect 29428 12684 29438 12740
rect 119200 12712 119800 12936
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 200 12040 800 12264
rect 101826 12012 101836 12068
rect 101892 12012 114940 12068
rect 114996 12012 115006 12068
rect 116274 11788 116284 11844
rect 116340 11788 116844 11844
rect 116900 11788 116910 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 116844 11620 116900 11788
rect 728 11592 1932 11620
rect 200 11564 1932 11592
rect 1988 11564 1998 11620
rect 116844 11592 119336 11620
rect 116844 11564 119800 11592
rect 200 11368 800 11564
rect 119200 11368 119800 11564
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 3042 10444 3052 10500
rect 3108 10444 3500 10500
rect 3556 10444 26124 10500
rect 26180 10444 26190 10500
rect 728 10248 1932 10276
rect 200 10220 1932 10248
rect 1988 10220 1998 10276
rect 200 10024 800 10220
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 119200 10024 119800 10248
rect 115490 9548 115500 9604
rect 115556 9576 119336 9604
rect 115556 9548 119800 9576
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 119200 9352 119800 9548
rect 15362 9212 15372 9268
rect 15428 9212 37772 9268
rect 37828 9212 37838 9268
rect 56354 9212 56364 9268
rect 56420 9212 100268 9268
rect 100324 9212 100334 9268
rect 200 8680 800 8904
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 200 8008 800 8232
rect 102452 8204 114492 8260
rect 114548 8204 114940 8260
rect 114996 8204 115006 8260
rect 115826 8204 115836 8260
rect 115892 8232 119336 8260
rect 115892 8204 119800 8232
rect 102452 8036 102508 8204
rect 64754 7980 64764 8036
rect 64820 7980 102508 8036
rect 119200 8008 119800 8204
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 728 6888 1820 6916
rect 200 6860 1820 6888
rect 1876 6860 1886 6916
rect 115490 6860 115500 6916
rect 115556 6888 119336 6916
rect 115556 6860 119800 6888
rect 200 6664 800 6860
rect 98242 6748 98252 6804
rect 98308 6748 114828 6804
rect 114884 6748 114894 6804
rect 43586 6636 43596 6692
rect 43652 6636 46060 6692
rect 46116 6636 46126 6692
rect 119200 6664 119800 6860
rect 3042 6412 3052 6468
rect 3108 6412 3612 6468
rect 3668 6412 29484 6468
rect 29540 6412 29550 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 116162 6188 116172 6244
rect 116228 6188 116732 6244
rect 116788 6216 119336 6244
rect 116788 6188 119800 6216
rect 59938 5964 59948 6020
rect 60004 5964 114940 6020
rect 114996 5964 115006 6020
rect 119200 5992 119800 6188
rect 3042 5852 3052 5908
rect 3108 5852 3500 5908
rect 3556 5852 17836 5908
rect 17892 5852 17902 5908
rect 83122 5852 83132 5908
rect 83188 5852 96348 5908
rect 96404 5852 96414 5908
rect 112354 5852 112364 5908
rect 112420 5852 113148 5908
rect 113204 5852 113214 5908
rect 3826 5740 3836 5796
rect 3892 5740 5180 5796
rect 5236 5740 5246 5796
rect 104962 5740 104972 5796
rect 105028 5740 115500 5796
rect 115556 5740 115566 5796
rect 728 5544 1932 5572
rect 200 5516 1932 5544
rect 1988 5516 1998 5572
rect 200 5320 800 5516
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 4946 5180 4956 5236
rect 5012 5180 6076 5236
rect 6132 5180 8428 5236
rect 28130 5180 28140 5236
rect 28196 5180 34524 5236
rect 34580 5180 34590 5236
rect 41570 5180 41580 5236
rect 41636 5180 43260 5236
rect 43316 5180 43326 5236
rect 48514 5180 48524 5236
rect 48580 5180 49196 5236
rect 49252 5180 49756 5236
rect 49812 5180 49822 5236
rect 8372 5124 8428 5180
rect 4834 5068 4844 5124
rect 4900 5068 5628 5124
rect 5684 5068 6524 5124
rect 6580 5068 6590 5124
rect 8372 5068 20972 5124
rect 21028 5068 21038 5124
rect 26338 5068 26348 5124
rect 26404 5068 26908 5124
rect 26964 5068 36092 5124
rect 36148 5068 36158 5124
rect 62738 5068 62748 5124
rect 62804 5068 63980 5124
rect 64036 5068 64046 5124
rect 42354 4956 42364 5012
rect 42420 4956 48076 5012
rect 48132 4956 48412 5012
rect 48468 4956 48478 5012
rect 54002 4956 54012 5012
rect 54068 4956 54796 5012
rect 54852 4956 55244 5012
rect 55300 4956 55468 5012
rect 99138 4956 99148 5012
rect 99204 4956 99932 5012
rect 99988 4956 99998 5012
rect 104290 4956 104300 5012
rect 104356 4956 111356 5012
rect 111412 4956 111916 5012
rect 111972 4956 114268 5012
rect 116274 4956 116284 5012
rect 116340 4956 117292 5012
rect 117348 4956 117358 5012
rect 55412 4900 55468 4956
rect 55412 4844 81676 4900
rect 81732 4844 81742 4900
rect 112242 4844 112252 4900
rect 112308 4844 113148 4900
rect 113204 4844 113214 4900
rect 114212 4788 114268 4956
rect 116162 4844 116172 4900
rect 116228 4844 117068 4900
rect 117124 4872 119336 4900
rect 117124 4844 119800 4872
rect 114212 4732 116844 4788
rect 116900 4732 117404 4788
rect 117460 4732 117470 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 119200 4648 119800 4844
rect 11218 4508 11228 4564
rect 11284 4508 11900 4564
rect 11956 4508 42028 4564
rect 42084 4508 42364 4564
rect 42420 4508 42430 4564
rect 49410 4508 49420 4564
rect 49476 4508 50316 4564
rect 50372 4508 51660 4564
rect 51716 4508 51726 4564
rect 59826 4508 59836 4564
rect 59892 4508 61068 4564
rect 61124 4508 61134 4564
rect 81666 4508 81676 4564
rect 81732 4508 83468 4564
rect 83524 4508 90524 4564
rect 90580 4508 90590 4564
rect 101378 4508 101388 4564
rect 101444 4508 101454 4564
rect 103282 4508 103292 4564
rect 103348 4508 114268 4564
rect 117282 4508 117292 4564
rect 117348 4508 118860 4564
rect 118916 4508 118926 4564
rect 802 4396 812 4452
rect 868 4396 1932 4452
rect 1988 4396 2380 4452
rect 2436 4396 2446 4452
rect 3378 4396 3388 4452
rect 3444 4396 14252 4452
rect 14308 4396 14318 4452
rect 59490 4396 59500 4452
rect 59556 4396 67788 4452
rect 67844 4396 67854 4452
rect 70578 4396 70588 4452
rect 70644 4396 71820 4452
rect 71876 4396 71886 4452
rect 86594 4396 86604 4452
rect 86660 4396 87948 4452
rect 88004 4396 88014 4452
rect 92642 4396 92652 4452
rect 92708 4396 93996 4452
rect 94052 4396 94062 4452
rect 98018 4396 98028 4452
rect 98084 4396 99372 4452
rect 99428 4396 99438 4452
rect 101388 4340 101444 4508
rect 114212 4452 114268 4508
rect 102452 4396 103516 4452
rect 103572 4396 104300 4452
rect 104356 4396 104366 4452
rect 114212 4396 114940 4452
rect 114996 4396 115006 4452
rect 116274 4396 116284 4452
rect 116340 4396 117852 4452
rect 117908 4396 117918 4452
rect 102452 4340 102508 4396
rect 2818 4284 2828 4340
rect 2884 4284 3164 4340
rect 3220 4284 11228 4340
rect 11284 4284 11294 4340
rect 56578 4284 56588 4340
rect 56644 4284 57372 4340
rect 57428 4284 57438 4340
rect 78306 4284 78316 4340
rect 78372 4284 78876 4340
rect 78932 4284 78942 4340
rect 90178 4284 90188 4340
rect 90244 4284 98364 4340
rect 98420 4284 98430 4340
rect 99922 4284 99932 4340
rect 99988 4284 100940 4340
rect 100996 4284 102508 4340
rect 112354 4284 112364 4340
rect 112420 4284 117068 4340
rect 117124 4284 117134 4340
rect 728 4200 1820 4228
rect 200 4172 1820 4200
rect 1876 4172 1886 4228
rect 2146 4172 2156 4228
rect 2212 4172 3948 4228
rect 4004 4172 4014 4228
rect 8194 4172 8204 4228
rect 8260 4172 8764 4228
rect 8820 4172 45948 4228
rect 46004 4172 46014 4228
rect 54562 4172 54572 4228
rect 54628 4172 55468 4228
rect 55524 4172 55534 4228
rect 72706 4172 72716 4228
rect 72772 4172 74060 4228
rect 74116 4172 74126 4228
rect 78754 4172 78764 4228
rect 78820 4172 79548 4228
rect 79604 4172 79614 4228
rect 111682 4172 111692 4228
rect 111748 4172 117628 4228
rect 117684 4172 117694 4228
rect 200 3976 800 4172
rect 36530 4060 36540 4116
rect 36596 4060 54460 4116
rect 54516 4060 54526 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 19618 3836 19628 3892
rect 19684 3836 21532 3892
rect 21588 3836 21598 3892
rect 8372 3724 12908 3780
rect 12964 3724 12974 3780
rect 20626 3724 20636 3780
rect 20692 3724 34412 3780
rect 34468 3724 34478 3780
rect 63858 3724 63868 3780
rect 63924 3724 66780 3780
rect 66836 3724 66846 3780
rect 8372 3668 8428 3724
rect 130 3612 140 3668
rect 196 3612 2044 3668
rect 2100 3612 2110 3668
rect 4946 3612 4956 3668
rect 5012 3612 8428 3668
rect 11442 3612 11452 3668
rect 11508 3612 12236 3668
rect 12292 3612 12302 3668
rect 16482 3612 16492 3668
rect 16548 3612 24332 3668
rect 24388 3612 24398 3668
rect 48514 3612 48524 3668
rect 48580 3612 49532 3668
rect 49588 3612 49598 3668
rect 59490 3612 59500 3668
rect 59556 3612 60508 3668
rect 60564 3612 60574 3668
rect 102946 3612 102956 3668
rect 103012 3612 104412 3668
rect 104468 3612 104478 3668
rect 108322 3612 108332 3668
rect 108388 3612 111580 3668
rect 111636 3612 111646 3668
rect 728 3528 3724 3556
rect 200 3500 3724 3528
rect 3780 3500 3790 3556
rect 88498 3500 88508 3556
rect 88564 3500 89964 3556
rect 90020 3500 90030 3556
rect 100258 3500 100268 3556
rect 100324 3500 102620 3556
rect 102676 3500 102686 3556
rect 112354 3500 112364 3556
rect 112420 3500 113820 3556
rect 113876 3500 113886 3556
rect 117842 3500 117852 3556
rect 117908 3528 119336 3556
rect 117908 3500 119800 3528
rect 200 3304 800 3500
rect 2034 3388 2044 3444
rect 2100 3388 2828 3444
rect 2884 3388 2894 3444
rect 3490 3388 3500 3444
rect 3556 3388 6412 3444
rect 6468 3388 6478 3444
rect 8866 3388 8876 3444
rect 8932 3388 9772 3444
rect 9828 3388 9838 3444
rect 20962 3388 20972 3444
rect 21028 3388 21196 3444
rect 21252 3388 21532 3444
rect 21588 3388 21598 3444
rect 24658 3388 24668 3444
rect 24724 3388 25452 3444
rect 25508 3388 25518 3444
rect 44258 3388 44268 3444
rect 44324 3388 45164 3444
rect 45220 3388 45230 3444
rect 55458 3388 55468 3444
rect 55524 3388 55804 3444
rect 55860 3388 56588 3444
rect 56644 3388 56654 3444
rect 63298 3388 63308 3444
rect 63364 3388 64092 3444
rect 64148 3388 64158 3444
rect 69122 3388 69132 3444
rect 69188 3388 70476 3444
rect 70532 3388 70542 3444
rect 74050 3388 74060 3444
rect 74116 3388 75068 3444
rect 75124 3388 75740 3444
rect 75796 3388 75806 3444
rect 83458 3388 83468 3444
rect 83524 3388 85148 3444
rect 85204 3388 85214 3444
rect 91298 3388 91308 3444
rect 91364 3388 92988 3444
rect 93044 3388 93054 3444
rect 96002 3388 96012 3444
rect 96068 3388 97356 3444
rect 97412 3388 97422 3444
rect 100930 3388 100940 3444
rect 100996 3388 101724 3444
rect 101780 3388 101790 3444
rect 110898 3388 110908 3444
rect 110964 3388 112588 3444
rect 112644 3388 112654 3444
rect 114258 3388 114268 3444
rect 114324 3388 116508 3444
rect 116564 3388 116574 3444
rect 75394 3276 75404 3332
rect 75460 3276 76300 3332
rect 76356 3276 76366 3332
rect 119200 3304 119800 3500
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 728 2184 3500 2212
rect 200 2156 3500 2184
rect 3556 2156 3566 2212
rect 118066 2156 118076 2212
rect 118132 2184 119336 2212
rect 118132 2156 119800 2184
rect 200 1960 800 2156
rect 119200 1960 119800 2156
rect 114482 1484 114492 1540
rect 114548 1512 119336 1540
rect 114548 1484 119800 1512
rect 119200 1288 119800 1484
rect 200 616 800 840
rect 119200 -56 119800 168
<< via3 >>
rect 4476 116788 4532 116844
rect 4580 116788 4636 116844
rect 4684 116788 4740 116844
rect 35196 116788 35252 116844
rect 35300 116788 35356 116844
rect 35404 116788 35460 116844
rect 65916 116788 65972 116844
rect 66020 116788 66076 116844
rect 66124 116788 66180 116844
rect 96636 116788 96692 116844
rect 96740 116788 96796 116844
rect 96844 116788 96900 116844
rect 19836 116004 19892 116060
rect 19940 116004 19996 116060
rect 20044 116004 20100 116060
rect 50556 116004 50612 116060
rect 50660 116004 50716 116060
rect 50764 116004 50820 116060
rect 81276 116004 81332 116060
rect 81380 116004 81436 116060
rect 81484 116004 81540 116060
rect 111996 116004 112052 116060
rect 112100 116004 112156 116060
rect 112204 116004 112260 116060
rect 4476 115220 4532 115276
rect 4580 115220 4636 115276
rect 4684 115220 4740 115276
rect 35196 115220 35252 115276
rect 35300 115220 35356 115276
rect 35404 115220 35460 115276
rect 65916 115220 65972 115276
rect 66020 115220 66076 115276
rect 66124 115220 66180 115276
rect 96636 115220 96692 115276
rect 96740 115220 96796 115276
rect 96844 115220 96900 115276
rect 19836 114436 19892 114492
rect 19940 114436 19996 114492
rect 20044 114436 20100 114492
rect 50556 114436 50612 114492
rect 50660 114436 50716 114492
rect 50764 114436 50820 114492
rect 81276 114436 81332 114492
rect 81380 114436 81436 114492
rect 81484 114436 81540 114492
rect 111996 114436 112052 114492
rect 112100 114436 112156 114492
rect 112204 114436 112260 114492
rect 4476 113652 4532 113708
rect 4580 113652 4636 113708
rect 4684 113652 4740 113708
rect 35196 113652 35252 113708
rect 35300 113652 35356 113708
rect 35404 113652 35460 113708
rect 65916 113652 65972 113708
rect 66020 113652 66076 113708
rect 66124 113652 66180 113708
rect 96636 113652 96692 113708
rect 96740 113652 96796 113708
rect 96844 113652 96900 113708
rect 19836 112868 19892 112924
rect 19940 112868 19996 112924
rect 20044 112868 20100 112924
rect 50556 112868 50612 112924
rect 50660 112868 50716 112924
rect 50764 112868 50820 112924
rect 81276 112868 81332 112924
rect 81380 112868 81436 112924
rect 81484 112868 81540 112924
rect 111996 112868 112052 112924
rect 112100 112868 112156 112924
rect 112204 112868 112260 112924
rect 4476 112084 4532 112140
rect 4580 112084 4636 112140
rect 4684 112084 4740 112140
rect 35196 112084 35252 112140
rect 35300 112084 35356 112140
rect 35404 112084 35460 112140
rect 65916 112084 65972 112140
rect 66020 112084 66076 112140
rect 66124 112084 66180 112140
rect 96636 112084 96692 112140
rect 96740 112084 96796 112140
rect 96844 112084 96900 112140
rect 19836 111300 19892 111356
rect 19940 111300 19996 111356
rect 20044 111300 20100 111356
rect 50556 111300 50612 111356
rect 50660 111300 50716 111356
rect 50764 111300 50820 111356
rect 81276 111300 81332 111356
rect 81380 111300 81436 111356
rect 81484 111300 81540 111356
rect 111996 111300 112052 111356
rect 112100 111300 112156 111356
rect 112204 111300 112260 111356
rect 4476 110516 4532 110572
rect 4580 110516 4636 110572
rect 4684 110516 4740 110572
rect 35196 110516 35252 110572
rect 35300 110516 35356 110572
rect 35404 110516 35460 110572
rect 65916 110516 65972 110572
rect 66020 110516 66076 110572
rect 66124 110516 66180 110572
rect 96636 110516 96692 110572
rect 96740 110516 96796 110572
rect 96844 110516 96900 110572
rect 19836 109732 19892 109788
rect 19940 109732 19996 109788
rect 20044 109732 20100 109788
rect 50556 109732 50612 109788
rect 50660 109732 50716 109788
rect 50764 109732 50820 109788
rect 81276 109732 81332 109788
rect 81380 109732 81436 109788
rect 81484 109732 81540 109788
rect 111996 109732 112052 109788
rect 112100 109732 112156 109788
rect 112204 109732 112260 109788
rect 4476 108948 4532 109004
rect 4580 108948 4636 109004
rect 4684 108948 4740 109004
rect 35196 108948 35252 109004
rect 35300 108948 35356 109004
rect 35404 108948 35460 109004
rect 65916 108948 65972 109004
rect 66020 108948 66076 109004
rect 66124 108948 66180 109004
rect 96636 108948 96692 109004
rect 96740 108948 96796 109004
rect 96844 108948 96900 109004
rect 19836 108164 19892 108220
rect 19940 108164 19996 108220
rect 20044 108164 20100 108220
rect 50556 108164 50612 108220
rect 50660 108164 50716 108220
rect 50764 108164 50820 108220
rect 81276 108164 81332 108220
rect 81380 108164 81436 108220
rect 81484 108164 81540 108220
rect 111996 108164 112052 108220
rect 112100 108164 112156 108220
rect 112204 108164 112260 108220
rect 4476 107380 4532 107436
rect 4580 107380 4636 107436
rect 4684 107380 4740 107436
rect 35196 107380 35252 107436
rect 35300 107380 35356 107436
rect 35404 107380 35460 107436
rect 65916 107380 65972 107436
rect 66020 107380 66076 107436
rect 66124 107380 66180 107436
rect 96636 107380 96692 107436
rect 96740 107380 96796 107436
rect 96844 107380 96900 107436
rect 19836 106596 19892 106652
rect 19940 106596 19996 106652
rect 20044 106596 20100 106652
rect 50556 106596 50612 106652
rect 50660 106596 50716 106652
rect 50764 106596 50820 106652
rect 81276 106596 81332 106652
rect 81380 106596 81436 106652
rect 81484 106596 81540 106652
rect 111996 106596 112052 106652
rect 112100 106596 112156 106652
rect 112204 106596 112260 106652
rect 4476 105812 4532 105868
rect 4580 105812 4636 105868
rect 4684 105812 4740 105868
rect 35196 105812 35252 105868
rect 35300 105812 35356 105868
rect 35404 105812 35460 105868
rect 65916 105812 65972 105868
rect 66020 105812 66076 105868
rect 66124 105812 66180 105868
rect 96636 105812 96692 105868
rect 96740 105812 96796 105868
rect 96844 105812 96900 105868
rect 19836 105028 19892 105084
rect 19940 105028 19996 105084
rect 20044 105028 20100 105084
rect 50556 105028 50612 105084
rect 50660 105028 50716 105084
rect 50764 105028 50820 105084
rect 81276 105028 81332 105084
rect 81380 105028 81436 105084
rect 81484 105028 81540 105084
rect 111996 105028 112052 105084
rect 112100 105028 112156 105084
rect 112204 105028 112260 105084
rect 4476 104244 4532 104300
rect 4580 104244 4636 104300
rect 4684 104244 4740 104300
rect 35196 104244 35252 104300
rect 35300 104244 35356 104300
rect 35404 104244 35460 104300
rect 65916 104244 65972 104300
rect 66020 104244 66076 104300
rect 66124 104244 66180 104300
rect 96636 104244 96692 104300
rect 96740 104244 96796 104300
rect 96844 104244 96900 104300
rect 19836 103460 19892 103516
rect 19940 103460 19996 103516
rect 20044 103460 20100 103516
rect 50556 103460 50612 103516
rect 50660 103460 50716 103516
rect 50764 103460 50820 103516
rect 81276 103460 81332 103516
rect 81380 103460 81436 103516
rect 81484 103460 81540 103516
rect 111996 103460 112052 103516
rect 112100 103460 112156 103516
rect 112204 103460 112260 103516
rect 4476 102676 4532 102732
rect 4580 102676 4636 102732
rect 4684 102676 4740 102732
rect 35196 102676 35252 102732
rect 35300 102676 35356 102732
rect 35404 102676 35460 102732
rect 65916 102676 65972 102732
rect 66020 102676 66076 102732
rect 66124 102676 66180 102732
rect 96636 102676 96692 102732
rect 96740 102676 96796 102732
rect 96844 102676 96900 102732
rect 19836 101892 19892 101948
rect 19940 101892 19996 101948
rect 20044 101892 20100 101948
rect 50556 101892 50612 101948
rect 50660 101892 50716 101948
rect 50764 101892 50820 101948
rect 81276 101892 81332 101948
rect 81380 101892 81436 101948
rect 81484 101892 81540 101948
rect 111996 101892 112052 101948
rect 112100 101892 112156 101948
rect 112204 101892 112260 101948
rect 4476 101108 4532 101164
rect 4580 101108 4636 101164
rect 4684 101108 4740 101164
rect 35196 101108 35252 101164
rect 35300 101108 35356 101164
rect 35404 101108 35460 101164
rect 65916 101108 65972 101164
rect 66020 101108 66076 101164
rect 66124 101108 66180 101164
rect 96636 101108 96692 101164
rect 96740 101108 96796 101164
rect 96844 101108 96900 101164
rect 19836 100324 19892 100380
rect 19940 100324 19996 100380
rect 20044 100324 20100 100380
rect 50556 100324 50612 100380
rect 50660 100324 50716 100380
rect 50764 100324 50820 100380
rect 81276 100324 81332 100380
rect 81380 100324 81436 100380
rect 81484 100324 81540 100380
rect 111996 100324 112052 100380
rect 112100 100324 112156 100380
rect 112204 100324 112260 100380
rect 4476 99540 4532 99596
rect 4580 99540 4636 99596
rect 4684 99540 4740 99596
rect 35196 99540 35252 99596
rect 35300 99540 35356 99596
rect 35404 99540 35460 99596
rect 65916 99540 65972 99596
rect 66020 99540 66076 99596
rect 66124 99540 66180 99596
rect 96636 99540 96692 99596
rect 96740 99540 96796 99596
rect 96844 99540 96900 99596
rect 19836 98756 19892 98812
rect 19940 98756 19996 98812
rect 20044 98756 20100 98812
rect 50556 98756 50612 98812
rect 50660 98756 50716 98812
rect 50764 98756 50820 98812
rect 81276 98756 81332 98812
rect 81380 98756 81436 98812
rect 81484 98756 81540 98812
rect 111996 98756 112052 98812
rect 112100 98756 112156 98812
rect 112204 98756 112260 98812
rect 4476 97972 4532 98028
rect 4580 97972 4636 98028
rect 4684 97972 4740 98028
rect 35196 97972 35252 98028
rect 35300 97972 35356 98028
rect 35404 97972 35460 98028
rect 65916 97972 65972 98028
rect 66020 97972 66076 98028
rect 66124 97972 66180 98028
rect 96636 97972 96692 98028
rect 96740 97972 96796 98028
rect 96844 97972 96900 98028
rect 19836 97188 19892 97244
rect 19940 97188 19996 97244
rect 20044 97188 20100 97244
rect 50556 97188 50612 97244
rect 50660 97188 50716 97244
rect 50764 97188 50820 97244
rect 81276 97188 81332 97244
rect 81380 97188 81436 97244
rect 81484 97188 81540 97244
rect 111996 97188 112052 97244
rect 112100 97188 112156 97244
rect 112204 97188 112260 97244
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 65916 96404 65972 96460
rect 66020 96404 66076 96460
rect 66124 96404 66180 96460
rect 96636 96404 96692 96460
rect 96740 96404 96796 96460
rect 96844 96404 96900 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 50556 95620 50612 95676
rect 50660 95620 50716 95676
rect 50764 95620 50820 95676
rect 81276 95620 81332 95676
rect 81380 95620 81436 95676
rect 81484 95620 81540 95676
rect 111996 95620 112052 95676
rect 112100 95620 112156 95676
rect 112204 95620 112260 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 65916 94836 65972 94892
rect 66020 94836 66076 94892
rect 66124 94836 66180 94892
rect 96636 94836 96692 94892
rect 96740 94836 96796 94892
rect 96844 94836 96900 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 50556 94052 50612 94108
rect 50660 94052 50716 94108
rect 50764 94052 50820 94108
rect 81276 94052 81332 94108
rect 81380 94052 81436 94108
rect 81484 94052 81540 94108
rect 111996 94052 112052 94108
rect 112100 94052 112156 94108
rect 112204 94052 112260 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 65916 93268 65972 93324
rect 66020 93268 66076 93324
rect 66124 93268 66180 93324
rect 96636 93268 96692 93324
rect 96740 93268 96796 93324
rect 96844 93268 96900 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 50556 92484 50612 92540
rect 50660 92484 50716 92540
rect 50764 92484 50820 92540
rect 81276 92484 81332 92540
rect 81380 92484 81436 92540
rect 81484 92484 81540 92540
rect 111996 92484 112052 92540
rect 112100 92484 112156 92540
rect 112204 92484 112260 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 65916 91700 65972 91756
rect 66020 91700 66076 91756
rect 66124 91700 66180 91756
rect 96636 91700 96692 91756
rect 96740 91700 96796 91756
rect 96844 91700 96900 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 50556 90916 50612 90972
rect 50660 90916 50716 90972
rect 50764 90916 50820 90972
rect 81276 90916 81332 90972
rect 81380 90916 81436 90972
rect 81484 90916 81540 90972
rect 111996 90916 112052 90972
rect 112100 90916 112156 90972
rect 112204 90916 112260 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 65916 90132 65972 90188
rect 66020 90132 66076 90188
rect 66124 90132 66180 90188
rect 96636 90132 96692 90188
rect 96740 90132 96796 90188
rect 96844 90132 96900 90188
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 50556 89348 50612 89404
rect 50660 89348 50716 89404
rect 50764 89348 50820 89404
rect 81276 89348 81332 89404
rect 81380 89348 81436 89404
rect 81484 89348 81540 89404
rect 111996 89348 112052 89404
rect 112100 89348 112156 89404
rect 112204 89348 112260 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 65916 88564 65972 88620
rect 66020 88564 66076 88620
rect 66124 88564 66180 88620
rect 96636 88564 96692 88620
rect 96740 88564 96796 88620
rect 96844 88564 96900 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 50556 87780 50612 87836
rect 50660 87780 50716 87836
rect 50764 87780 50820 87836
rect 81276 87780 81332 87836
rect 81380 87780 81436 87836
rect 81484 87780 81540 87836
rect 111996 87780 112052 87836
rect 112100 87780 112156 87836
rect 112204 87780 112260 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 65916 86996 65972 87052
rect 66020 86996 66076 87052
rect 66124 86996 66180 87052
rect 96636 86996 96692 87052
rect 96740 86996 96796 87052
rect 96844 86996 96900 87052
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 50556 86212 50612 86268
rect 50660 86212 50716 86268
rect 50764 86212 50820 86268
rect 81276 86212 81332 86268
rect 81380 86212 81436 86268
rect 81484 86212 81540 86268
rect 111996 86212 112052 86268
rect 112100 86212 112156 86268
rect 112204 86212 112260 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 65916 85428 65972 85484
rect 66020 85428 66076 85484
rect 66124 85428 66180 85484
rect 96636 85428 96692 85484
rect 96740 85428 96796 85484
rect 96844 85428 96900 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 50556 84644 50612 84700
rect 50660 84644 50716 84700
rect 50764 84644 50820 84700
rect 81276 84644 81332 84700
rect 81380 84644 81436 84700
rect 81484 84644 81540 84700
rect 111996 84644 112052 84700
rect 112100 84644 112156 84700
rect 112204 84644 112260 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 65916 83860 65972 83916
rect 66020 83860 66076 83916
rect 66124 83860 66180 83916
rect 96636 83860 96692 83916
rect 96740 83860 96796 83916
rect 96844 83860 96900 83916
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 50556 83076 50612 83132
rect 50660 83076 50716 83132
rect 50764 83076 50820 83132
rect 81276 83076 81332 83132
rect 81380 83076 81436 83132
rect 81484 83076 81540 83132
rect 111996 83076 112052 83132
rect 112100 83076 112156 83132
rect 112204 83076 112260 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 65916 82292 65972 82348
rect 66020 82292 66076 82348
rect 66124 82292 66180 82348
rect 96636 82292 96692 82348
rect 96740 82292 96796 82348
rect 96844 82292 96900 82348
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 50556 81508 50612 81564
rect 50660 81508 50716 81564
rect 50764 81508 50820 81564
rect 81276 81508 81332 81564
rect 81380 81508 81436 81564
rect 81484 81508 81540 81564
rect 111996 81508 112052 81564
rect 112100 81508 112156 81564
rect 112204 81508 112260 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 65916 80724 65972 80780
rect 66020 80724 66076 80780
rect 66124 80724 66180 80780
rect 96636 80724 96692 80780
rect 96740 80724 96796 80780
rect 96844 80724 96900 80780
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 50556 79940 50612 79996
rect 50660 79940 50716 79996
rect 50764 79940 50820 79996
rect 81276 79940 81332 79996
rect 81380 79940 81436 79996
rect 81484 79940 81540 79996
rect 111996 79940 112052 79996
rect 112100 79940 112156 79996
rect 112204 79940 112260 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 65916 79156 65972 79212
rect 66020 79156 66076 79212
rect 66124 79156 66180 79212
rect 96636 79156 96692 79212
rect 96740 79156 96796 79212
rect 96844 79156 96900 79212
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 50556 78372 50612 78428
rect 50660 78372 50716 78428
rect 50764 78372 50820 78428
rect 81276 78372 81332 78428
rect 81380 78372 81436 78428
rect 81484 78372 81540 78428
rect 111996 78372 112052 78428
rect 112100 78372 112156 78428
rect 112204 78372 112260 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 65916 77588 65972 77644
rect 66020 77588 66076 77644
rect 66124 77588 66180 77644
rect 96636 77588 96692 77644
rect 96740 77588 96796 77644
rect 96844 77588 96900 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 81276 76804 81332 76860
rect 81380 76804 81436 76860
rect 81484 76804 81540 76860
rect 111996 76804 112052 76860
rect 112100 76804 112156 76860
rect 112204 76804 112260 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 96636 76020 96692 76076
rect 96740 76020 96796 76076
rect 96844 76020 96900 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 81276 75236 81332 75292
rect 81380 75236 81436 75292
rect 81484 75236 81540 75292
rect 111996 75236 112052 75292
rect 112100 75236 112156 75292
rect 112204 75236 112260 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 96636 74452 96692 74508
rect 96740 74452 96796 74508
rect 96844 74452 96900 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 81276 73668 81332 73724
rect 81380 73668 81436 73724
rect 81484 73668 81540 73724
rect 111996 73668 112052 73724
rect 112100 73668 112156 73724
rect 112204 73668 112260 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 96636 72884 96692 72940
rect 96740 72884 96796 72940
rect 96844 72884 96900 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 81276 72100 81332 72156
rect 81380 72100 81436 72156
rect 81484 72100 81540 72156
rect 111996 72100 112052 72156
rect 112100 72100 112156 72156
rect 112204 72100 112260 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 96636 71316 96692 71372
rect 96740 71316 96796 71372
rect 96844 71316 96900 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 81276 70532 81332 70588
rect 81380 70532 81436 70588
rect 81484 70532 81540 70588
rect 111996 70532 112052 70588
rect 112100 70532 112156 70588
rect 112204 70532 112260 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 96636 69748 96692 69804
rect 96740 69748 96796 69804
rect 96844 69748 96900 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 81276 68964 81332 69020
rect 81380 68964 81436 69020
rect 81484 68964 81540 69020
rect 111996 68964 112052 69020
rect 112100 68964 112156 69020
rect 112204 68964 112260 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 96636 68180 96692 68236
rect 96740 68180 96796 68236
rect 96844 68180 96900 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 81276 67396 81332 67452
rect 81380 67396 81436 67452
rect 81484 67396 81540 67452
rect 111996 67396 112052 67452
rect 112100 67396 112156 67452
rect 112204 67396 112260 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 96636 66612 96692 66668
rect 96740 66612 96796 66668
rect 96844 66612 96900 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 81276 65828 81332 65884
rect 81380 65828 81436 65884
rect 81484 65828 81540 65884
rect 111996 65828 112052 65884
rect 112100 65828 112156 65884
rect 112204 65828 112260 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 96636 65044 96692 65100
rect 96740 65044 96796 65100
rect 96844 65044 96900 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 81276 64260 81332 64316
rect 81380 64260 81436 64316
rect 81484 64260 81540 64316
rect 111996 64260 112052 64316
rect 112100 64260 112156 64316
rect 112204 64260 112260 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 96636 63476 96692 63532
rect 96740 63476 96796 63532
rect 96844 63476 96900 63532
rect 73276 63308 73332 63364
rect 73276 63084 73332 63140
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 81276 62692 81332 62748
rect 81380 62692 81436 62748
rect 81484 62692 81540 62748
rect 111996 62692 112052 62748
rect 112100 62692 112156 62748
rect 112204 62692 112260 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 96636 61908 96692 61964
rect 96740 61908 96796 61964
rect 96844 61908 96900 61964
rect 59388 61628 59444 61684
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 81276 61124 81332 61180
rect 81380 61124 81436 61180
rect 81484 61124 81540 61180
rect 111996 61124 112052 61180
rect 112100 61124 112156 61180
rect 112204 61124 112260 61180
rect 55468 60620 55524 60676
rect 58492 60508 58548 60564
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 96636 60340 96692 60396
rect 96740 60340 96796 60396
rect 96844 60340 96900 60396
rect 55468 60284 55524 60340
rect 59388 59948 59444 60004
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 81276 59556 81332 59612
rect 81380 59556 81436 59612
rect 81484 59556 81540 59612
rect 111996 59556 112052 59612
rect 112100 59556 112156 59612
rect 112204 59556 112260 59612
rect 58492 59388 58548 59444
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 96636 58772 96692 58828
rect 96740 58772 96796 58828
rect 96844 58772 96900 58828
rect 62524 58604 62580 58660
rect 62076 58492 62132 58548
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 81276 57988 81332 58044
rect 81380 57988 81436 58044
rect 81484 57988 81540 58044
rect 111996 57988 112052 58044
rect 112100 57988 112156 58044
rect 112204 57988 112260 58044
rect 49868 57820 49924 57876
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 96636 57204 96692 57260
rect 96740 57204 96796 57260
rect 96844 57204 96900 57260
rect 51212 57148 51268 57204
rect 65100 56812 65156 56868
rect 49980 56588 50036 56644
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 111996 56420 112052 56476
rect 112100 56420 112156 56476
rect 112204 56420 112260 56476
rect 65100 55916 65156 55972
rect 50988 55804 51044 55860
rect 51100 55692 51156 55748
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 50316 55580 50372 55636
rect 55132 55468 55188 55524
rect 62748 55132 62804 55188
rect 50204 55020 50260 55076
rect 51212 55020 51268 55076
rect 50988 54908 51044 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 111996 54852 112052 54908
rect 112100 54852 112156 54908
rect 112204 54852 112260 54908
rect 51772 54796 51828 54852
rect 55132 54796 55188 54852
rect 58492 54796 58548 54852
rect 62748 54796 62804 54852
rect 49868 54460 49924 54516
rect 50316 54460 50372 54516
rect 51100 54460 51156 54516
rect 50204 54236 50260 54292
rect 51212 54236 51268 54292
rect 51772 54236 51828 54292
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 62412 53676 62468 53732
rect 58492 53452 58548 53508
rect 62412 53340 62468 53396
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 111996 53284 112052 53340
rect 112100 53284 112156 53340
rect 112204 53284 112260 53340
rect 49980 52892 50036 52948
rect 53228 52780 53284 52836
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 47740 52108 47796 52164
rect 49980 51884 50036 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 111996 51716 112052 51772
rect 112100 51716 112156 51772
rect 112204 51716 112260 51772
rect 52444 51100 52500 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 55916 50876 55972 50932
rect 61852 50764 61908 50820
rect 65100 50764 65156 50820
rect 51212 50540 51268 50596
rect 61852 50428 61908 50484
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 111996 50148 112052 50204
rect 112100 50148 112156 50204
rect 112204 50148 112260 50204
rect 52556 49980 52612 50036
rect 52556 49644 52612 49700
rect 53228 49420 53284 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 60844 49196 60900 49252
rect 67452 48972 67508 49028
rect 60844 48748 60900 48804
rect 52444 48636 52500 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 111996 48580 112052 48636
rect 112100 48580 112156 48636
rect 112204 48580 112260 48636
rect 67452 48524 67508 48580
rect 57148 48412 57204 48468
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 55916 47404 55972 47460
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 111996 47012 112052 47068
rect 112100 47012 112156 47068
rect 112204 47012 112260 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 47740 46172 47796 46228
rect 51212 45500 51268 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 57148 45276 57204 45332
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 62188 44044 62244 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 62076 43708 62132 43764
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
<< metal4 >>
rect 4448 116844 4768 116876
rect 4448 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4768 116844
rect 4448 115276 4768 116788
rect 4448 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4768 115276
rect 4448 113708 4768 115220
rect 4448 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4768 113708
rect 4448 112140 4768 113652
rect 4448 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4768 112140
rect 4448 110572 4768 112084
rect 4448 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4768 110572
rect 4448 109004 4768 110516
rect 4448 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4768 109004
rect 4448 107436 4768 108948
rect 4448 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4768 107436
rect 4448 105868 4768 107380
rect 4448 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4768 105868
rect 4448 104300 4768 105812
rect 4448 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4768 104300
rect 4448 102732 4768 104244
rect 4448 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4768 102732
rect 4448 101164 4768 102676
rect 4448 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4768 101164
rect 4448 99596 4768 101108
rect 4448 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4768 99596
rect 4448 98028 4768 99540
rect 4448 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4768 98028
rect 4448 96460 4768 97972
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 116060 20128 116876
rect 19808 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20128 116060
rect 19808 114492 20128 116004
rect 19808 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20128 114492
rect 19808 112924 20128 114436
rect 19808 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20128 112924
rect 19808 111356 20128 112868
rect 19808 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20128 111356
rect 19808 109788 20128 111300
rect 19808 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20128 109788
rect 19808 108220 20128 109732
rect 19808 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20128 108220
rect 19808 106652 20128 108164
rect 19808 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20128 106652
rect 19808 105084 20128 106596
rect 19808 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20128 105084
rect 19808 103516 20128 105028
rect 19808 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20128 103516
rect 19808 101948 20128 103460
rect 19808 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20128 101948
rect 19808 100380 20128 101892
rect 19808 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20128 100380
rect 19808 98812 20128 100324
rect 19808 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20128 98812
rect 19808 97244 20128 98756
rect 19808 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20128 97244
rect 19808 95676 20128 97188
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 116844 35488 116876
rect 35168 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35488 116844
rect 35168 115276 35488 116788
rect 35168 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35488 115276
rect 35168 113708 35488 115220
rect 35168 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35488 113708
rect 35168 112140 35488 113652
rect 35168 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35488 112140
rect 35168 110572 35488 112084
rect 35168 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35488 110572
rect 35168 109004 35488 110516
rect 35168 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35488 109004
rect 35168 107436 35488 108948
rect 35168 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35488 107436
rect 35168 105868 35488 107380
rect 35168 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35488 105868
rect 35168 104300 35488 105812
rect 35168 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35488 104300
rect 35168 102732 35488 104244
rect 35168 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35488 102732
rect 35168 101164 35488 102676
rect 35168 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35488 101164
rect 35168 99596 35488 101108
rect 35168 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35488 99596
rect 35168 98028 35488 99540
rect 35168 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35488 98028
rect 35168 96460 35488 97972
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 50528 116060 50848 116876
rect 50528 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50848 116060
rect 50528 114492 50848 116004
rect 50528 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50848 114492
rect 50528 112924 50848 114436
rect 50528 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50848 112924
rect 50528 111356 50848 112868
rect 50528 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50848 111356
rect 50528 109788 50848 111300
rect 50528 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50848 109788
rect 50528 108220 50848 109732
rect 50528 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50848 108220
rect 50528 106652 50848 108164
rect 50528 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50848 106652
rect 50528 105084 50848 106596
rect 50528 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50848 105084
rect 50528 103516 50848 105028
rect 50528 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50848 103516
rect 50528 101948 50848 103460
rect 50528 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50848 101948
rect 50528 100380 50848 101892
rect 50528 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50848 100380
rect 50528 98812 50848 100324
rect 50528 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50848 98812
rect 50528 97244 50848 98756
rect 50528 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50848 97244
rect 50528 95676 50848 97188
rect 50528 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50848 95676
rect 50528 94108 50848 95620
rect 50528 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50848 94108
rect 50528 92540 50848 94052
rect 50528 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50848 92540
rect 50528 90972 50848 92484
rect 50528 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50848 90972
rect 50528 89404 50848 90916
rect 50528 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50848 89404
rect 50528 87836 50848 89348
rect 50528 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50848 87836
rect 50528 86268 50848 87780
rect 50528 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50848 86268
rect 50528 84700 50848 86212
rect 50528 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50848 84700
rect 50528 83132 50848 84644
rect 50528 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50848 83132
rect 50528 81564 50848 83076
rect 50528 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50848 81564
rect 50528 79996 50848 81508
rect 50528 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50848 79996
rect 50528 78428 50848 79940
rect 50528 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50848 78428
rect 50528 76860 50848 78372
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 65888 116844 66208 116876
rect 65888 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66208 116844
rect 65888 115276 66208 116788
rect 65888 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66208 115276
rect 65888 113708 66208 115220
rect 65888 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66208 113708
rect 65888 112140 66208 113652
rect 65888 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66208 112140
rect 65888 110572 66208 112084
rect 65888 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66208 110572
rect 65888 109004 66208 110516
rect 65888 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66208 109004
rect 65888 107436 66208 108948
rect 65888 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66208 107436
rect 65888 105868 66208 107380
rect 65888 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66208 105868
rect 65888 104300 66208 105812
rect 65888 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66208 104300
rect 65888 102732 66208 104244
rect 65888 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66208 102732
rect 65888 101164 66208 102676
rect 65888 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66208 101164
rect 65888 99596 66208 101108
rect 65888 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66208 99596
rect 65888 98028 66208 99540
rect 65888 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66208 98028
rect 65888 96460 66208 97972
rect 65888 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66208 96460
rect 65888 94892 66208 96404
rect 65888 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66208 94892
rect 65888 93324 66208 94836
rect 65888 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66208 93324
rect 65888 91756 66208 93268
rect 65888 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66208 91756
rect 65888 90188 66208 91700
rect 65888 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66208 90188
rect 65888 88620 66208 90132
rect 65888 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66208 88620
rect 65888 87052 66208 88564
rect 65888 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66208 87052
rect 65888 85484 66208 86996
rect 65888 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66208 85484
rect 65888 83916 66208 85428
rect 65888 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66208 83916
rect 65888 82348 66208 83860
rect 65888 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66208 82348
rect 65888 80780 66208 82292
rect 65888 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66208 80780
rect 65888 79212 66208 80724
rect 65888 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66208 79212
rect 65888 77644 66208 79156
rect 65888 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66208 77644
rect 65888 76076 66208 77588
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 81248 116060 81568 116876
rect 81248 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81568 116060
rect 81248 114492 81568 116004
rect 81248 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81568 114492
rect 81248 112924 81568 114436
rect 81248 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81568 112924
rect 81248 111356 81568 112868
rect 81248 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81568 111356
rect 81248 109788 81568 111300
rect 81248 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81568 109788
rect 81248 108220 81568 109732
rect 81248 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81568 108220
rect 81248 106652 81568 108164
rect 81248 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81568 106652
rect 81248 105084 81568 106596
rect 81248 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81568 105084
rect 81248 103516 81568 105028
rect 81248 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81568 103516
rect 81248 101948 81568 103460
rect 81248 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81568 101948
rect 81248 100380 81568 101892
rect 81248 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81568 100380
rect 81248 98812 81568 100324
rect 81248 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81568 98812
rect 81248 97244 81568 98756
rect 81248 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81568 97244
rect 81248 95676 81568 97188
rect 81248 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81568 95676
rect 81248 94108 81568 95620
rect 81248 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81568 94108
rect 81248 92540 81568 94052
rect 81248 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81568 92540
rect 81248 90972 81568 92484
rect 81248 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81568 90972
rect 81248 89404 81568 90916
rect 81248 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81568 89404
rect 81248 87836 81568 89348
rect 81248 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81568 87836
rect 81248 86268 81568 87780
rect 81248 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81568 86268
rect 81248 84700 81568 86212
rect 81248 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81568 84700
rect 81248 83132 81568 84644
rect 81248 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81568 83132
rect 81248 81564 81568 83076
rect 81248 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81568 81564
rect 81248 79996 81568 81508
rect 81248 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81568 79996
rect 81248 78428 81568 79940
rect 81248 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81568 78428
rect 81248 76860 81568 78372
rect 81248 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81568 76860
rect 81248 75292 81568 76804
rect 81248 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81568 75292
rect 81248 73724 81568 75236
rect 81248 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81568 73724
rect 81248 72156 81568 73668
rect 81248 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81568 72156
rect 81248 70588 81568 72100
rect 81248 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81568 70588
rect 81248 69020 81568 70532
rect 81248 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81568 69020
rect 81248 67452 81568 68964
rect 81248 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81568 67452
rect 81248 65884 81568 67396
rect 81248 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81568 65884
rect 81248 64316 81568 65828
rect 81248 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81568 64316
rect 73276 63364 73332 63374
rect 73276 63140 73332 63308
rect 73276 63074 73332 63084
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 59388 61684 59444 61694
rect 55468 60676 55524 60686
rect 55468 60340 55524 60620
rect 55468 60274 55524 60284
rect 58492 60564 58548 60574
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 58492 59444 58548 60508
rect 59388 60004 59444 61628
rect 59388 59938 59444 59948
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 58492 59378 58548 59388
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 62524 58660 62580 58670
rect 62076 58548 62132 58558
rect 62524 58548 62580 58604
rect 62132 58492 62580 58548
rect 62076 58482 62132 58492
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 49868 57876 49924 57886
rect 49868 54516 49924 57820
rect 49868 54450 49924 54460
rect 49980 56644 50036 56654
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 49980 52948 50036 56588
rect 50528 56476 50848 57988
rect 65888 57260 66208 58772
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50316 55636 50372 55646
rect 50204 55076 50260 55086
rect 50204 54292 50260 55020
rect 50316 54516 50372 55580
rect 50316 54450 50372 54460
rect 50528 54908 50848 56420
rect 51212 57204 51268 57214
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50988 55860 51044 55870
rect 50988 54964 51044 55804
rect 50988 54898 51044 54908
rect 51100 55748 51156 55758
rect 50204 54226 50260 54236
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 47740 52164 47796 52174
rect 47740 46228 47796 52108
rect 49980 51940 50036 52892
rect 49980 51874 50036 51884
rect 50528 53340 50848 54852
rect 51100 54516 51156 55692
rect 51100 54450 51156 54460
rect 51212 55076 51268 57148
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65100 56868 65156 56878
rect 65100 55972 65156 56812
rect 51212 54292 51268 55020
rect 55132 55524 55188 55534
rect 51212 54226 51268 54236
rect 51772 54852 51828 54862
rect 51772 54292 51828 54796
rect 55132 54852 55188 55468
rect 62748 55188 62804 55198
rect 55132 54786 55188 54796
rect 58492 54852 58548 54862
rect 51772 54226 51828 54236
rect 58492 53508 58548 54796
rect 62748 54852 62804 55132
rect 62748 54786 62804 54796
rect 58492 53442 58548 53452
rect 62412 53732 62468 53742
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 62412 53396 62468 53676
rect 62412 53330 62468 53340
rect 47740 46162 47796 46172
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 53228 52836 53284 52846
rect 52444 51156 52500 51166
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 51212 50596 51268 50606
rect 51212 45556 51268 50540
rect 52444 48692 52500 51100
rect 52556 50036 52612 50046
rect 52556 49700 52612 49980
rect 52556 49634 52612 49644
rect 53228 49476 53284 52780
rect 53228 49410 53284 49420
rect 55916 50932 55972 50942
rect 52444 48626 52500 48636
rect 55916 47460 55972 50876
rect 61852 50820 61908 50830
rect 61852 50484 61908 50764
rect 65100 50820 65156 55916
rect 65100 50754 65156 50764
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 61852 50418 61908 50428
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 60844 49252 60900 49262
rect 60844 48804 60900 49196
rect 60844 48738 60900 48748
rect 55916 47394 55972 47404
rect 57148 48468 57204 48478
rect 51212 45490 51268 45500
rect 50528 43932 50848 45444
rect 57148 45332 57204 48412
rect 57148 45266 57204 45276
rect 65888 47852 66208 49364
rect 81248 62748 81568 64260
rect 81248 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81568 62748
rect 81248 61180 81568 62692
rect 81248 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81568 61180
rect 81248 59612 81568 61124
rect 81248 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81568 59612
rect 81248 58044 81568 59556
rect 81248 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81568 58044
rect 81248 56476 81568 57988
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 67452 49028 67508 49038
rect 67452 48580 67508 48972
rect 67452 48514 67508 48524
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 62188 44100 62244 44110
rect 62076 43764 62132 43774
rect 62188 43764 62244 44044
rect 62132 43708 62244 43764
rect 62076 43698 62132 43708
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 47068 81568 48580
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 116844 96928 116876
rect 96608 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96928 116844
rect 96608 115276 96928 116788
rect 96608 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96928 115276
rect 96608 113708 96928 115220
rect 96608 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96928 113708
rect 96608 112140 96928 113652
rect 96608 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96928 112140
rect 96608 110572 96928 112084
rect 96608 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96928 110572
rect 96608 109004 96928 110516
rect 96608 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96928 109004
rect 96608 107436 96928 108948
rect 96608 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96928 107436
rect 96608 105868 96928 107380
rect 96608 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96928 105868
rect 96608 104300 96928 105812
rect 96608 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96928 104300
rect 96608 102732 96928 104244
rect 96608 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96928 102732
rect 96608 101164 96928 102676
rect 96608 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96928 101164
rect 96608 99596 96928 101108
rect 96608 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96928 99596
rect 96608 98028 96928 99540
rect 96608 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96928 98028
rect 96608 96460 96928 97972
rect 96608 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96928 96460
rect 96608 94892 96928 96404
rect 96608 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96928 94892
rect 96608 93324 96928 94836
rect 96608 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96928 93324
rect 96608 91756 96928 93268
rect 96608 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96928 91756
rect 96608 90188 96928 91700
rect 96608 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96928 90188
rect 96608 88620 96928 90132
rect 96608 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96928 88620
rect 96608 87052 96928 88564
rect 96608 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96928 87052
rect 96608 85484 96928 86996
rect 96608 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96928 85484
rect 96608 83916 96928 85428
rect 96608 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96928 83916
rect 96608 82348 96928 83860
rect 96608 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96928 82348
rect 96608 80780 96928 82292
rect 96608 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96928 80780
rect 96608 79212 96928 80724
rect 96608 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96928 79212
rect 96608 77644 96928 79156
rect 96608 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96928 77644
rect 96608 76076 96928 77588
rect 96608 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96928 76076
rect 96608 74508 96928 76020
rect 96608 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96928 74508
rect 96608 72940 96928 74452
rect 96608 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96928 72940
rect 96608 71372 96928 72884
rect 96608 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96928 71372
rect 96608 69804 96928 71316
rect 96608 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96928 69804
rect 96608 68236 96928 69748
rect 96608 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96928 68236
rect 96608 66668 96928 68180
rect 96608 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96928 66668
rect 96608 65100 96928 66612
rect 96608 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96928 65100
rect 96608 63532 96928 65044
rect 96608 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96928 63532
rect 96608 61964 96928 63476
rect 96608 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96928 61964
rect 96608 60396 96928 61908
rect 96608 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96928 60396
rect 96608 58828 96928 60340
rect 96608 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96928 58828
rect 96608 57260 96928 58772
rect 96608 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96928 57260
rect 96608 55692 96928 57204
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 96608 54124 96928 55636
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 111968 116060 112288 116876
rect 111968 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112288 116060
rect 111968 114492 112288 116004
rect 111968 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112288 114492
rect 111968 112924 112288 114436
rect 111968 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112288 112924
rect 111968 111356 112288 112868
rect 111968 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112288 111356
rect 111968 109788 112288 111300
rect 111968 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112288 109788
rect 111968 108220 112288 109732
rect 111968 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112288 108220
rect 111968 106652 112288 108164
rect 111968 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112288 106652
rect 111968 105084 112288 106596
rect 111968 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112288 105084
rect 111968 103516 112288 105028
rect 111968 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112288 103516
rect 111968 101948 112288 103460
rect 111968 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112288 101948
rect 111968 100380 112288 101892
rect 111968 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112288 100380
rect 111968 98812 112288 100324
rect 111968 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112288 98812
rect 111968 97244 112288 98756
rect 111968 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112288 97244
rect 111968 95676 112288 97188
rect 111968 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112288 95676
rect 111968 94108 112288 95620
rect 111968 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112288 94108
rect 111968 92540 112288 94052
rect 111968 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112288 92540
rect 111968 90972 112288 92484
rect 111968 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112288 90972
rect 111968 89404 112288 90916
rect 111968 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112288 89404
rect 111968 87836 112288 89348
rect 111968 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112288 87836
rect 111968 86268 112288 87780
rect 111968 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112288 86268
rect 111968 84700 112288 86212
rect 111968 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112288 84700
rect 111968 83132 112288 84644
rect 111968 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112288 83132
rect 111968 81564 112288 83076
rect 111968 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112288 81564
rect 111968 79996 112288 81508
rect 111968 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112288 79996
rect 111968 78428 112288 79940
rect 111968 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112288 78428
rect 111968 76860 112288 78372
rect 111968 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112288 76860
rect 111968 75292 112288 76804
rect 111968 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112288 75292
rect 111968 73724 112288 75236
rect 111968 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112288 73724
rect 111968 72156 112288 73668
rect 111968 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112288 72156
rect 111968 70588 112288 72100
rect 111968 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112288 70588
rect 111968 69020 112288 70532
rect 111968 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112288 69020
rect 111968 67452 112288 68964
rect 111968 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112288 67452
rect 111968 65884 112288 67396
rect 111968 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112288 65884
rect 111968 64316 112288 65828
rect 111968 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112288 64316
rect 111968 62748 112288 64260
rect 111968 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112288 62748
rect 111968 61180 112288 62692
rect 111968 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112288 61180
rect 111968 59612 112288 61124
rect 111968 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112288 59612
rect 111968 58044 112288 59556
rect 111968 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112288 58044
rect 111968 56476 112288 57988
rect 111968 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112288 56476
rect 111968 54908 112288 56420
rect 111968 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112288 54908
rect 111968 53340 112288 54852
rect 111968 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112288 53340
rect 111968 51772 112288 53284
rect 111968 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112288 51772
rect 111968 50204 112288 51716
rect 111968 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112288 50204
rect 111968 48636 112288 50148
rect 111968 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112288 48636
rect 111968 47068 112288 48580
rect 111968 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112288 47068
rect 111968 45500 112288 47012
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 111968 11004 112288 12516
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 111968 4732 112288 6244
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 111968 3164 112288 4676
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__I gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 67200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1669390400
transform 1 0 65744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A1
timestamp 1669390400
transform -1 0 37968 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A2
timestamp 1669390400
transform -1 0 39536 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1669390400
transform 1 0 41104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1669390400
transform 1 0 51408 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1669390400
transform -1 0 51968 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A2
timestamp 1669390400
transform 1 0 63168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1669390400
transform 1 0 60928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__I
timestamp 1669390400
transform 1 0 49280 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1669390400
transform 1 0 70560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1669390400
transform 1 0 45472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__I
timestamp 1669390400
transform 1 0 48272 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A1
timestamp 1669390400
transform 1 0 45024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A2
timestamp 1669390400
transform -1 0 46144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A1
timestamp 1669390400
transform -1 0 45584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A2
timestamp 1669390400
transform -1 0 45136 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I0
timestamp 1669390400
transform 1 0 93072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I1
timestamp 1669390400
transform 1 0 90496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__S
timestamp 1669390400
transform 1 0 90048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__I1
timestamp 1669390400
transform 1 0 115360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__S
timestamp 1669390400
transform 1 0 114912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I0
timestamp 1669390400
transform -1 0 45584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I1
timestamp 1669390400
transform 1 0 47712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__S
timestamp 1669390400
transform 1 0 48160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I0
timestamp 1669390400
transform -1 0 45584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I1
timestamp 1669390400
transform 1 0 47712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__S
timestamp 1669390400
transform -1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1669390400
transform 1 0 49392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I0
timestamp 1669390400
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I1
timestamp 1669390400
transform 1 0 47376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__S
timestamp 1669390400
transform 1 0 47824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I0
timestamp 1669390400
transform 1 0 117824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I1
timestamp 1669390400
transform 1 0 114352 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__S
timestamp 1669390400
transform 1 0 113456 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__I
timestamp 1669390400
transform 1 0 70112 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A1
timestamp 1669390400
transform 1 0 73248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A2
timestamp 1669390400
transform -1 0 71904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A1
timestamp 1669390400
transform -1 0 69664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A2
timestamp 1669390400
transform 1 0 71008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__I0
timestamp 1669390400
transform 1 0 79520 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__I1
timestamp 1669390400
transform 1 0 77168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__S
timestamp 1669390400
transform 1 0 77392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__I0
timestamp 1669390400
transform 1 0 76496 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__I1
timestamp 1669390400
transform 1 0 74144 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__S
timestamp 1669390400
transform 1 0 74592 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__I
timestamp 1669390400
transform 1 0 66304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A1
timestamp 1669390400
transform -1 0 68768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A2
timestamp 1669390400
transform 1 0 68096 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A2
timestamp 1669390400
transform 1 0 68432 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I0
timestamp 1669390400
transform 1 0 47376 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I1
timestamp 1669390400
transform -1 0 47152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__S
timestamp 1669390400
transform 1 0 46480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__I0
timestamp 1669390400
transform 1 0 115472 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__I1
timestamp 1669390400
transform 1 0 115920 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__S
timestamp 1669390400
transform -1 0 117152 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__I0
timestamp 1669390400
transform 1 0 73248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__I1
timestamp 1669390400
transform 1 0 70672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__S
timestamp 1669390400
transform 1 0 70224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__I
timestamp 1669390400
transform 1 0 49952 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A1
timestamp 1669390400
transform 1 0 73696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A2
timestamp 1669390400
transform 1 0 73248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A1
timestamp 1669390400
transform -1 0 70560 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A2
timestamp 1669390400
transform 1 0 72688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__I
timestamp 1669390400
transform 1 0 67312 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A1
timestamp 1669390400
transform 1 0 72128 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A2
timestamp 1669390400
transform 1 0 71232 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A1
timestamp 1669390400
transform 1 0 69440 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A2
timestamp 1669390400
transform 1 0 71680 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I0
timestamp 1669390400
transform 1 0 45360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I1
timestamp 1669390400
transform 1 0 47712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__S
timestamp 1669390400
transform 1 0 48160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I0
timestamp 1669390400
transform -1 0 56112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I1
timestamp 1669390400
transform 1 0 56336 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__S
timestamp 1669390400
transform 1 0 53536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I0
timestamp 1669390400
transform 1 0 80192 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I1
timestamp 1669390400
transform 1 0 77840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__S
timestamp 1669390400
transform 1 0 78288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I0
timestamp 1669390400
transform 1 0 44688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I1
timestamp 1669390400
transform 1 0 47376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__S
timestamp 1669390400
transform 1 0 47824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I0
timestamp 1669390400
transform -1 0 45808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I1
timestamp 1669390400
transform -1 0 45920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__S
timestamp 1669390400
transform 1 0 47824 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I0
timestamp 1669390400
transform 1 0 44688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I1
timestamp 1669390400
transform 1 0 47264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__S
timestamp 1669390400
transform 1 0 47936 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1669390400
transform 1 0 49168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1669390400
transform 1 0 49616 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A2
timestamp 1669390400
transform 1 0 49168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1669390400
transform -1 0 50736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A2
timestamp 1669390400
transform -1 0 48832 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__I
timestamp 1669390400
transform -1 0 52528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A1
timestamp 1669390400
transform 1 0 45696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A2
timestamp 1669390400
transform -1 0 46368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A2
timestamp 1669390400
transform 1 0 45248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__I0
timestamp 1669390400
transform 1 0 47376 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__I1
timestamp 1669390400
transform -1 0 49952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__S
timestamp 1669390400
transform 1 0 50176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__I
timestamp 1669390400
transform -1 0 48496 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__A1
timestamp 1669390400
transform 1 0 46928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__A2
timestamp 1669390400
transform 1 0 48048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A2
timestamp 1669390400
transform -1 0 46928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__I0
timestamp 1669390400
transform 1 0 64064 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__I1
timestamp 1669390400
transform 1 0 60592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__S
timestamp 1669390400
transform -1 0 63168 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__I0
timestamp 1669390400
transform 1 0 49616 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__I1
timestamp 1669390400
transform -1 0 49392 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__S
timestamp 1669390400
transform 1 0 51296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I0
timestamp 1669390400
transform 1 0 63840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I1
timestamp 1669390400
transform 1 0 61040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__S
timestamp 1669390400
transform 1 0 63392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__I
timestamp 1669390400
transform 1 0 71344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A1
timestamp 1669390400
transform -1 0 74368 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A2
timestamp 1669390400
transform 1 0 73024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A2
timestamp 1669390400
transform 1 0 71792 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__I
timestamp 1669390400
transform 1 0 68880 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__A1
timestamp 1669390400
transform 1 0 51184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__A2
timestamp 1669390400
transform -1 0 50288 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A1
timestamp 1669390400
transform 1 0 51072 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A2
timestamp 1669390400
transform 1 0 49504 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__I
timestamp 1669390400
transform 1 0 70896 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1669390400
transform -1 0 74816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A2
timestamp 1669390400
transform 1 0 74144 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__A2
timestamp 1669390400
transform 1 0 71008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A1
timestamp 1669390400
transform 1 0 52752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2
timestamp 1669390400
transform 1 0 56112 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__A1
timestamp 1669390400
transform 1 0 53648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__A2
timestamp 1669390400
transform -1 0 49728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1669390400
transform -1 0 69888 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A2
timestamp 1669390400
transform 1 0 69216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__A1
timestamp 1669390400
transform 1 0 65296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__A2
timestamp 1669390400
transform -1 0 64288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1669390400
transform -1 0 67312 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A2
timestamp 1669390400
transform 1 0 66864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__I
timestamp 1669390400
transform 1 0 61488 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__A2
timestamp 1669390400
transform 1 0 60368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A1
timestamp 1669390400
transform -1 0 53536 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A2
timestamp 1669390400
transform 1 0 52640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A1
timestamp 1669390400
transform 1 0 56448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1669390400
transform -1 0 53312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A2
timestamp 1669390400
transform -1 0 52080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A1
timestamp 1669390400
transform -1 0 55664 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A2
timestamp 1669390400
transform 1 0 54992 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1
timestamp 1669390400
transform 1 0 52192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1669390400
transform -1 0 53760 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A1
timestamp 1669390400
transform 1 0 40320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A2
timestamp 1669390400
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A1
timestamp 1669390400
transform -1 0 39760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A2
timestamp 1669390400
transform 1 0 39984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A1
timestamp 1669390400
transform -1 0 71008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A2
timestamp 1669390400
transform 1 0 69216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A1
timestamp 1669390400
transform 1 0 48272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A2
timestamp 1669390400
transform 1 0 50960 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__B
timestamp 1669390400
transform 1 0 48160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A1
timestamp 1669390400
transform -1 0 52416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A2
timestamp 1669390400
transform -1 0 49280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A3
timestamp 1669390400
transform -1 0 50624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A1
timestamp 1669390400
transform -1 0 50960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A2
timestamp 1669390400
transform 1 0 51184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A3
timestamp 1669390400
transform -1 0 51968 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__A1
timestamp 1669390400
transform 1 0 62048 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__A2
timestamp 1669390400
transform 1 0 61600 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A1
timestamp 1669390400
transform -1 0 64624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A2
timestamp 1669390400
transform 1 0 61600 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1669390400
transform -1 0 58128 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1669390400
transform -1 0 59024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1669390400
transform 1 0 52192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A2
timestamp 1669390400
transform 1 0 52640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A1
timestamp 1669390400
transform 1 0 61264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A2
timestamp 1669390400
transform 1 0 60480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A4
timestamp 1669390400
transform 1 0 59696 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A1
timestamp 1669390400
transform -1 0 62832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A2
timestamp 1669390400
transform 1 0 62160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A1
timestamp 1669390400
transform -1 0 69552 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A2
timestamp 1669390400
transform -1 0 68320 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A1
timestamp 1669390400
transform 1 0 62384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A2
timestamp 1669390400
transform 1 0 61936 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A1
timestamp 1669390400
transform 1 0 57568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A2
timestamp 1669390400
transform 1 0 59472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A1
timestamp 1669390400
transform 1 0 63952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A2
timestamp 1669390400
transform -1 0 63280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A3
timestamp 1669390400
transform 1 0 60592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__A1
timestamp 1669390400
transform 1 0 60032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__A2
timestamp 1669390400
transform 1 0 60480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A1
timestamp 1669390400
transform 1 0 42000 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A2
timestamp 1669390400
transform 1 0 42448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__A1
timestamp 1669390400
transform -1 0 64288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__A2
timestamp 1669390400
transform 1 0 64288 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A1
timestamp 1669390400
transform -1 0 57792 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A2
timestamp 1669390400
transform -1 0 56000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A2
timestamp 1669390400
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A4
timestamp 1669390400
transform 1 0 60032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1669390400
transform -1 0 59024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A2
timestamp 1669390400
transform 1 0 60368 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__B
timestamp 1669390400
transform 1 0 59248 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1669390400
transform -1 0 60816 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A2
timestamp 1669390400
transform 1 0 60032 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A1
timestamp 1669390400
transform -1 0 58688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A2
timestamp 1669390400
transform 1 0 54656 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__B
timestamp 1669390400
transform 1 0 55552 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1669390400
transform -1 0 58576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1669390400
transform 1 0 56672 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__B
timestamp 1669390400
transform 1 0 60704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A2
timestamp 1669390400
transform -1 0 57680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A1
timestamp 1669390400
transform -1 0 52864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A1
timestamp 1669390400
transform 1 0 56896 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A2
timestamp 1669390400
transform 1 0 54992 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__B
timestamp 1669390400
transform 1 0 54544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__A1
timestamp 1669390400
transform -1 0 60592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__B1
timestamp 1669390400
transform -1 0 53872 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__B2
timestamp 1669390400
transform 1 0 62272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A1
timestamp 1669390400
transform -1 0 66864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A2
timestamp 1669390400
transform 1 0 65296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A3
timestamp 1669390400
transform -1 0 64624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1669390400
transform 1 0 55328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A2
timestamp 1669390400
transform 1 0 55888 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A1
timestamp 1669390400
transform 1 0 54432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A2
timestamp 1669390400
transform -1 0 54432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A3
timestamp 1669390400
transform -1 0 53760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A1
timestamp 1669390400
transform -1 0 56784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__B1
timestamp 1669390400
transform 1 0 54880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A1
timestamp 1669390400
transform -1 0 54208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__A1
timestamp 1669390400
transform 1 0 64512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__A2
timestamp 1669390400
transform 1 0 66640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__A1
timestamp 1669390400
transform 1 0 69216 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__A1
timestamp 1669390400
transform 1 0 65296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__B1
timestamp 1669390400
transform 1 0 67424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A1
timestamp 1669390400
transform -1 0 67872 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A2
timestamp 1669390400
transform 1 0 66192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A3
timestamp 1669390400
transform 1 0 65632 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A1
timestamp 1669390400
transform 1 0 65296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A2
timestamp 1669390400
transform 1 0 57568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A3
timestamp 1669390400
transform 1 0 61936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A1
timestamp 1669390400
transform 1 0 60928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A1
timestamp 1669390400
transform -1 0 57456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A2
timestamp 1669390400
transform -1 0 58352 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A3
timestamp 1669390400
transform 1 0 54656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A1
timestamp 1669390400
transform -1 0 56448 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A2
timestamp 1669390400
transform -1 0 56896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__B1
timestamp 1669390400
transform 1 0 55104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A1
timestamp 1669390400
transform 1 0 59584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1669390400
transform -1 0 58128 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A2
timestamp 1669390400
transform -1 0 58576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A1
timestamp 1669390400
transform -1 0 57680 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A1
timestamp 1669390400
transform 1 0 65296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1669390400
transform 1 0 64400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A3
timestamp 1669390400
transform 1 0 63504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A4
timestamp 1669390400
transform 1 0 63952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__A1
timestamp 1669390400
transform 1 0 57344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A1
timestamp 1669390400
transform 1 0 57680 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A2
timestamp 1669390400
transform -1 0 57568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A1
timestamp 1669390400
transform -1 0 56896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__B1
timestamp 1669390400
transform -1 0 58800 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__B2
timestamp 1669390400
transform 1 0 57120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A1
timestamp 1669390400
transform -1 0 57344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__B
timestamp 1669390400
transform 1 0 57456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__A1
timestamp 1669390400
transform 1 0 59024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A1
timestamp 1669390400
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A1
timestamp 1669390400
transform 1 0 58128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__B1
timestamp 1669390400
transform 1 0 56672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__C1
timestamp 1669390400
transform -1 0 56448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__C2
timestamp 1669390400
transform 1 0 60368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__A1
timestamp 1669390400
transform 1 0 63504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A1
timestamp 1669390400
transform -1 0 56000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1669390400
transform -1 0 54208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1669390400
transform 1 0 63056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1669390400
transform 1 0 60032 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A1
timestamp 1669390400
transform -1 0 64624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1669390400
transform -1 0 67312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A2
timestamp 1669390400
transform 1 0 66192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__B2
timestamp 1669390400
transform 1 0 60480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__B
timestamp 1669390400
transform 1 0 65744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__A1
timestamp 1669390400
transform 1 0 64848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__A2
timestamp 1669390400
transform 1 0 65296 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A1
timestamp 1669390400
transform -1 0 66304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A2
timestamp 1669390400
transform 1 0 66080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A3
timestamp 1669390400
transform 1 0 62160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A1
timestamp 1669390400
transform 1 0 64624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A2
timestamp 1669390400
transform 1 0 65744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A1
timestamp 1669390400
transform 1 0 62608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__B1
timestamp 1669390400
transform 1 0 62384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__C1
timestamp 1669390400
transform 1 0 62832 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__C2
timestamp 1669390400
transform -1 0 65520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1669390400
transform 1 0 65520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A1
timestamp 1669390400
transform -1 0 52528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A2
timestamp 1669390400
transform -1 0 52080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A1
timestamp 1669390400
transform 1 0 57904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1669390400
transform 1 0 56000 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A1
timestamp 1669390400
transform 1 0 66640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A2
timestamp 1669390400
transform 1 0 66192 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A1
timestamp 1669390400
transform 1 0 64288 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1669390400
transform -1 0 55328 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__A1
timestamp 1669390400
transform 1 0 65744 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__A2
timestamp 1669390400
transform -1 0 62944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__B1
timestamp 1669390400
transform 1 0 62272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__C1
timestamp 1669390400
transform 1 0 61824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__C2
timestamp 1669390400
transform -1 0 66864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A1
timestamp 1669390400
transform 1 0 65296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__A1
timestamp 1669390400
transform 1 0 64400 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__B
timestamp 1669390400
transform 1 0 64624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A1
timestamp 1669390400
transform 1 0 66528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A2
timestamp 1669390400
transform 1 0 67088 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__A1
timestamp 1669390400
transform -1 0 64848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__A2
timestamp 1669390400
transform -1 0 66304 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A1
timestamp 1669390400
transform 1 0 61376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A1
timestamp 1669390400
transform 1 0 59248 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__B1
timestamp 1669390400
transform 1 0 57680 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__B2
timestamp 1669390400
transform 1 0 60256 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__B
timestamp 1669390400
transform 1 0 62384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__A1
timestamp 1669390400
transform 1 0 64624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A1
timestamp 1669390400
transform 1 0 64512 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A2
timestamp 1669390400
transform 1 0 63840 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__B1
timestamp 1669390400
transform 1 0 62160 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__C1
timestamp 1669390400
transform 1 0 60928 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__C2
timestamp 1669390400
transform -1 0 61600 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A1
timestamp 1669390400
transform -1 0 64064 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__A2
timestamp 1669390400
transform 1 0 68432 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__A3
timestamp 1669390400
transform 1 0 68992 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__A1
timestamp 1669390400
transform 1 0 55664 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__A2
timestamp 1669390400
transform -1 0 55440 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A1
timestamp 1669390400
transform 1 0 56336 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A2
timestamp 1669390400
transform -1 0 53424 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__B1
timestamp 1669390400
transform 1 0 55888 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__C1
timestamp 1669390400
transform 1 0 56784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__C2
timestamp 1669390400
transform -1 0 52976 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A1
timestamp 1669390400
transform 1 0 53424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A1
timestamp 1669390400
transform 1 0 56560 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A2
timestamp 1669390400
transform -1 0 57568 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A1
timestamp 1669390400
transform 1 0 55888 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A1
timestamp 1669390400
transform 1 0 59360 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A2
timestamp 1669390400
transform -1 0 53872 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__B1
timestamp 1669390400
transform -1 0 54768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__C1
timestamp 1669390400
transform 1 0 54992 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__C2
timestamp 1669390400
transform -1 0 53424 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__A1
timestamp 1669390400
transform 1 0 54208 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A1
timestamp 1669390400
transform 1 0 56448 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A1
timestamp 1669390400
transform 1 0 57792 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A1
timestamp 1669390400
transform -1 0 54320 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A2
timestamp 1669390400
transform 1 0 58464 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__B1
timestamp 1669390400
transform 1 0 58016 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__C1
timestamp 1669390400
transform -1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__C2
timestamp 1669390400
transform -1 0 55776 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A1
timestamp 1669390400
transform 1 0 58912 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A1
timestamp 1669390400
transform 1 0 60144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A2
timestamp 1669390400
transform -1 0 54992 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A3
timestamp 1669390400
transform 1 0 60592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A4
timestamp 1669390400
transform -1 0 59920 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A1
timestamp 1669390400
transform -1 0 52304 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A2
timestamp 1669390400
transform -1 0 52864 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1669390400
transform -1 0 54432 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__B1
timestamp 1669390400
transform -1 0 56896 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__B2
timestamp 1669390400
transform 1 0 52192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__I
timestamp 1669390400
transform -1 0 53648 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A1
timestamp 1669390400
transform -1 0 53648 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A3
timestamp 1669390400
transform 1 0 52976 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A1
timestamp 1669390400
transform -1 0 52416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A2
timestamp 1669390400
transform -1 0 52864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A1
timestamp 1669390400
transform -1 0 52752 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A1
timestamp 1669390400
transform 1 0 58912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1669390400
transform 1 0 56672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__B1
timestamp 1669390400
transform 1 0 57344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__C1
timestamp 1669390400
transform 1 0 56672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__C2
timestamp 1669390400
transform 1 0 59584 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A1
timestamp 1669390400
transform 1 0 57568 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A1
timestamp 1669390400
transform -1 0 57344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A2
timestamp 1669390400
transform 1 0 59360 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A1
timestamp 1669390400
transform -1 0 61712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A2
timestamp 1669390400
transform -1 0 60256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A1
timestamp 1669390400
transform 1 0 63056 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A1
timestamp 1669390400
transform 1 0 56672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__A1
timestamp 1669390400
transform -1 0 57568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A1
timestamp 1669390400
transform 1 0 61712 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1669390400
transform -1 0 60704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A1
timestamp 1669390400
transform -1 0 53312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__B1
timestamp 1669390400
transform 1 0 61824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__C1
timestamp 1669390400
transform 1 0 58128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__C2
timestamp 1669390400
transform 1 0 61376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A1
timestamp 1669390400
transform 1 0 60480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__I
timestamp 1669390400
transform 1 0 51296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__A1
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__B
timestamp 1669390400
transform -1 0 52976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A1
timestamp 1669390400
transform 1 0 56672 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A2
timestamp 1669390400
transform 1 0 55776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A1
timestamp 1669390400
transform 1 0 61936 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A2
timestamp 1669390400
transform 1 0 56224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A3
timestamp 1669390400
transform 1 0 62832 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A3
timestamp 1669390400
transform 1 0 51408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A1
timestamp 1669390400
transform -1 0 51184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__B1
timestamp 1669390400
transform 1 0 51856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__B2
timestamp 1669390400
transform -1 0 53984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A1
timestamp 1669390400
transform -1 0 56896 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A1
timestamp 1669390400
transform 1 0 61264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A2
timestamp 1669390400
transform 1 0 60144 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A1
timestamp 1669390400
transform 1 0 61264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__B1
timestamp 1669390400
transform 1 0 63504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__C1
timestamp 1669390400
transform 1 0 60592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__C2
timestamp 1669390400
transform 1 0 65072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__A1
timestamp 1669390400
transform 1 0 64400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A1
timestamp 1669390400
transform -1 0 47376 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A2
timestamp 1669390400
transform 1 0 47600 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A3
timestamp 1669390400
transform -1 0 52752 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A1
timestamp 1669390400
transform 1 0 48608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A2
timestamp 1669390400
transform -1 0 48944 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__B
timestamp 1669390400
transform 1 0 50512 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__A2
timestamp 1669390400
transform -1 0 48496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__A1
timestamp 1669390400
transform -1 0 48496 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__A2
timestamp 1669390400
transform -1 0 48048 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__B1
timestamp 1669390400
transform -1 0 48944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__B2
timestamp 1669390400
transform 1 0 47376 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__A1
timestamp 1669390400
transform 1 0 47824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A1
timestamp 1669390400
transform 1 0 49952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A2
timestamp 1669390400
transform 1 0 52640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__A1
timestamp 1669390400
transform 1 0 48720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__A2
timestamp 1669390400
transform -1 0 52416 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__B1
timestamp 1669390400
transform -1 0 54208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__C1
timestamp 1669390400
transform -1 0 53760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__C2
timestamp 1669390400
transform -1 0 47824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__A1
timestamp 1669390400
transform 1 0 55664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A1
timestamp 1669390400
transform 1 0 50848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A2
timestamp 1669390400
transform 1 0 50400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1669390400
transform 1 0 48160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A2
timestamp 1669390400
transform 1 0 48608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A1
timestamp 1669390400
transform 1 0 53536 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A2
timestamp 1669390400
transform 1 0 49168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A3
timestamp 1669390400
transform 1 0 53200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A1
timestamp 1669390400
transform 1 0 54880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B
timestamp 1669390400
transform 1 0 52864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__C
timestamp 1669390400
transform 1 0 51296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__A1
timestamp 1669390400
transform -1 0 68544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__A2
timestamp 1669390400
transform 1 0 67872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B1
timestamp 1669390400
transform 1 0 66416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B2
timestamp 1669390400
transform -1 0 68320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A2
timestamp 1669390400
transform -1 0 56000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__B
timestamp 1669390400
transform 1 0 55328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__A1
timestamp 1669390400
transform 1 0 49056 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__A2
timestamp 1669390400
transform 1 0 49504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__A1
timestamp 1669390400
transform 1 0 48272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__A2
timestamp 1669390400
transform -1 0 48944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__B1
timestamp 1669390400
transform -1 0 48272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__C1
timestamp 1669390400
transform -1 0 51632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__C2
timestamp 1669390400
transform 1 0 48272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A1
timestamp 1669390400
transform -1 0 51408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A1
timestamp 1669390400
transform 1 0 67872 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A2
timestamp 1669390400
transform 1 0 67424 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1669390400
transform -1 0 46144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A2
timestamp 1669390400
transform -1 0 47040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__A1
timestamp 1669390400
transform 1 0 69664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__A2
timestamp 1669390400
transform 1 0 67536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A1
timestamp 1669390400
transform -1 0 68320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__B1
timestamp 1669390400
transform 1 0 66416 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__C1
timestamp 1669390400
transform 1 0 65968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__C2
timestamp 1669390400
transform -1 0 67424 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A1
timestamp 1669390400
transform 1 0 67312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__A1
timestamp 1669390400
transform 1 0 52640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__A2
timestamp 1669390400
transform 1 0 49504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__A1
timestamp 1669390400
transform -1 0 51632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__A1
timestamp 1669390400
transform -1 0 56672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__A1
timestamp 1669390400
transform 1 0 68096 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__A2
timestamp 1669390400
transform 1 0 68544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__A1
timestamp 1669390400
transform 1 0 68544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A1
timestamp 1669390400
transform 1 0 57344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__A1
timestamp 1669390400
transform 1 0 68320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__B1
timestamp 1669390400
transform -1 0 67312 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__C1
timestamp 1669390400
transform 1 0 68320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__C2
timestamp 1669390400
transform 1 0 69664 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A1
timestamp 1669390400
transform 1 0 70112 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A1
timestamp 1669390400
transform -1 0 46592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A2
timestamp 1669390400
transform 1 0 48720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A1
timestamp 1669390400
transform -1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A2
timestamp 1669390400
transform -1 0 48496 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A3
timestamp 1669390400
transform -1 0 48944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__I
timestamp 1669390400
transform -1 0 49840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A1
timestamp 1669390400
transform 1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A2
timestamp 1669390400
transform 1 0 49168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A1
timestamp 1669390400
transform 1 0 48720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A3
timestamp 1669390400
transform 1 0 52640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__C
timestamp 1669390400
transform 1 0 47376 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__A1
timestamp 1669390400
transform -1 0 46480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B1
timestamp 1669390400
transform 1 0 47824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B2
timestamp 1669390400
transform 1 0 51520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A1
timestamp 1669390400
transform 1 0 46928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A1
timestamp 1669390400
transform 1 0 50960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A2
timestamp 1669390400
transform -1 0 51632 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A1
timestamp 1669390400
transform -1 0 48048 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A2
timestamp 1669390400
transform 1 0 48272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__B1
timestamp 1669390400
transform -1 0 50960 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__C1
timestamp 1669390400
transform 1 0 48720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__C2
timestamp 1669390400
transform 1 0 51184 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1669390400
transform 1 0 48720 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__A1
timestamp 1669390400
transform -1 0 46032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__A2
timestamp 1669390400
transform -1 0 46256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__A3
timestamp 1669390400
transform 1 0 47264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A1
timestamp 1669390400
transform 1 0 47376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A2
timestamp 1669390400
transform -1 0 47152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__B
timestamp 1669390400
transform 1 0 46480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__I
timestamp 1669390400
transform -1 0 70000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A1
timestamp 1669390400
transform 1 0 68544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A3
timestamp 1669390400
transform 1 0 66528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__A1
timestamp 1669390400
transform 1 0 45360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__A2
timestamp 1669390400
transform -1 0 46480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__C
timestamp 1669390400
transform -1 0 46928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A1
timestamp 1669390400
transform -1 0 47040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__A1
timestamp 1669390400
transform -1 0 48944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__A2
timestamp 1669390400
transform -1 0 48496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__A1
timestamp 1669390400
transform 1 0 47712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__A1
timestamp 1669390400
transform 1 0 46032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__B1
timestamp 1669390400
transform -1 0 50288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__C1
timestamp 1669390400
transform 1 0 46480 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__C2
timestamp 1669390400
transform -1 0 45808 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__579__A1
timestamp 1669390400
transform 1 0 50512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A1
timestamp 1669390400
transform 1 0 67200 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A2
timestamp 1669390400
transform 1 0 67648 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A3
timestamp 1669390400
transform 1 0 68096 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A4
timestamp 1669390400
transform 1 0 69216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A1
timestamp 1669390400
transform 1 0 71904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__A1
timestamp 1669390400
transform 1 0 71456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__A2
timestamp 1669390400
transform 1 0 71008 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__B1
timestamp 1669390400
transform 1 0 69104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__C1
timestamp 1669390400
transform 1 0 68656 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__C2
timestamp 1669390400
transform 1 0 71904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A1
timestamp 1669390400
transform 1 0 71232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A1
timestamp 1669390400
transform 1 0 71120 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A2
timestamp 1669390400
transform 1 0 71568 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A1
timestamp 1669390400
transform 1 0 70896 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A2
timestamp 1669390400
transform 1 0 68544 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A3
timestamp 1669390400
transform 1 0 68432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A4
timestamp 1669390400
transform 1 0 70560 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__B
timestamp 1669390400
transform 1 0 70448 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A1
timestamp 1669390400
transform 1 0 71680 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A1
timestamp 1669390400
transform -1 0 67872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A2
timestamp 1669390400
transform 1 0 71008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__B1
timestamp 1669390400
transform 1 0 68544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__B2
timestamp 1669390400
transform 1 0 71456 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__B
timestamp 1669390400
transform 1 0 68544 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A1
timestamp 1669390400
transform 1 0 71008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A2
timestamp 1669390400
transform 1 0 71456 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A3
timestamp 1669390400
transform -1 0 72128 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A2
timestamp 1669390400
transform 1 0 70448 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__A1
timestamp 1669390400
transform 1 0 67984 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__A1
timestamp 1669390400
transform 1 0 66192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__A2
timestamp 1669390400
transform 1 0 67088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A1
timestamp 1669390400
transform 1 0 70000 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__B1
timestamp 1669390400
transform 1 0 66976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__B2
timestamp 1669390400
transform 1 0 68320 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__B
timestamp 1669390400
transform 1 0 67536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__CLK
timestamp 1669390400
transform 1 0 70560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__D
timestamp 1669390400
transform 1 0 73696 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__CLK
timestamp 1669390400
transform 1 0 45808 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__CLK
timestamp 1669390400
transform 1 0 90608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__CLK
timestamp 1669390400
transform 1 0 114576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__CLK
timestamp 1669390400
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__CLK
timestamp 1669390400
transform -1 0 49056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__CLK
timestamp 1669390400
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__CLK
timestamp 1669390400
transform 1 0 113904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__CLK
timestamp 1669390400
transform 1 0 68992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__CLK
timestamp 1669390400
transform 1 0 81200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__CLK
timestamp 1669390400
transform -1 0 78400 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__607__CLK
timestamp 1669390400
transform 1 0 65296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__CLK
timestamp 1669390400
transform 1 0 48832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__CLK
timestamp 1669390400
transform 1 0 113904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__CLK
timestamp 1669390400
transform 1 0 75040 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__CLK
timestamp 1669390400
transform -1 0 74144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__CLK
timestamp 1669390400
transform 1 0 69216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__613__CLK
timestamp 1669390400
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__CLK
timestamp 1669390400
transform -1 0 52864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__CLK
timestamp 1669390400
transform 1 0 76496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__CLK
timestamp 1669390400
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__CLK
timestamp 1669390400
transform 1 0 46928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__CLK
timestamp 1669390400
transform -1 0 50064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__CLK
timestamp 1669390400
transform -1 0 49616 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__CLK
timestamp 1669390400
transform 1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__CLK
timestamp 1669390400
transform 1 0 49392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__CLK
timestamp 1669390400
transform 1 0 49392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__CLK
timestamp 1669390400
transform 1 0 64512 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__CLK
timestamp 1669390400
transform 1 0 50624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__CLK
timestamp 1669390400
transform 1 0 60592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__626__CLK
timestamp 1669390400
transform 1 0 74928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__CLK
timestamp 1669390400
transform 1 0 51968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__CLK
timestamp 1669390400
transform 1 0 74928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__CLK
timestamp 1669390400
transform 1 0 65184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__630__CLK
timestamp 1669390400
transform 1 0 54208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__CLK
timestamp 1669390400
transform -1 0 68096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__CLK
timestamp 1669390400
transform 1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__CLK
timestamp 1669390400
transform -1 0 62832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__CLK
timestamp 1669390400
transform 1 0 60592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__CLK
timestamp 1669390400
transform 1 0 67536 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__CLK
timestamp 1669390400
transform -1 0 66304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__637__CLK
timestamp 1669390400
transform 1 0 63056 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__CLK
timestamp 1669390400
transform 1 0 63056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__CLK
timestamp 1669390400
transform 1 0 66752 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__CLK
timestamp 1669390400
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__641__CLK
timestamp 1669390400
transform -1 0 55328 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__CLK
timestamp 1669390400
transform 1 0 60592 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__CLK
timestamp 1669390400
transform 1 0 51296 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__CLK
timestamp 1669390400
transform 1 0 62160 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__CLK
timestamp 1669390400
transform -1 0 65520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__CLK
timestamp 1669390400
transform 1 0 52640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__CLK
timestamp 1669390400
transform 1 0 62608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__648__CLK
timestamp 1669390400
transform 1 0 50512 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__CLK
timestamp 1669390400
transform 1 0 53312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__CLK
timestamp 1669390400
transform 1 0 53088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__CLK
timestamp 1669390400
transform 1 0 54432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__CLK
timestamp 1669390400
transform 1 0 69216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__CLK
timestamp 1669390400
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__CLK
timestamp 1669390400
transform 1 0 50960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__CLK
timestamp 1669390400
transform 1 0 50960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__CLK
timestamp 1669390400
transform 1 0 46368 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__CLK
timestamp 1669390400
transform 1 0 51408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__CLK
timestamp 1669390400
transform 1 0 73248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__CLK
timestamp 1669390400
transform 1 0 73472 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__660__CLK
timestamp 1669390400
transform 1 0 67984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__I
timestamp 1669390400
transform 1 0 4368 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__I
timestamp 1669390400
transform 1 0 116704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__I
timestamp 1669390400
transform -1 0 76608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__I
timestamp 1669390400
transform 1 0 116928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__I
timestamp 1669390400
transform 1 0 5264 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__I
timestamp 1669390400
transform 1 0 117040 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__I
timestamp 1669390400
transform 1 0 56896 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__I
timestamp 1669390400
transform 1 0 116816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__I
timestamp 1669390400
transform 1 0 116928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__I
timestamp 1669390400
transform 1 0 116256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__I
timestamp 1669390400
transform 1 0 3248 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__I
timestamp 1669390400
transform 1 0 3248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__I
timestamp 1669390400
transform 1 0 3248 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__I
timestamp 1669390400
transform 1 0 104272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__I
timestamp 1669390400
transform 1 0 117376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__I
timestamp 1669390400
transform 1 0 64064 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__I
timestamp 1669390400
transform -1 0 3472 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__I
timestamp 1669390400
transform 1 0 9744 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__I
timestamp 1669390400
transform 1 0 3248 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__I
timestamp 1669390400
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__I
timestamp 1669390400
transform 1 0 101360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__I
timestamp 1669390400
transform 1 0 11872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__I
timestamp 1669390400
transform 1 0 116256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__I
timestamp 1669390400
transform 1 0 3248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__I
timestamp 1669390400
transform 1 0 116704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__I
timestamp 1669390400
transform 1 0 42000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__I
timestamp 1669390400
transform 1 0 99904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__I
timestamp 1669390400
transform 1 0 3248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__I
timestamp 1669390400
transform 1 0 3248 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__I
timestamp 1669390400
transform 1 0 23744 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__I
timestamp 1669390400
transform -1 0 2128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__I
timestamp 1669390400
transform 1 0 116704 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__I
timestamp 1669390400
transform 1 0 116704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__I
timestamp 1669390400
transform 1 0 3248 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__I
timestamp 1669390400
transform 1 0 3248 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__I
timestamp 1669390400
transform 1 0 66304 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__I
timestamp 1669390400
transform 1 0 111328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__I
timestamp 1669390400
transform 1 0 34384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__741__I
timestamp 1669390400
transform 1 0 55216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__I
timestamp 1669390400
transform -1 0 116704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__I
timestamp 1669390400
transform -1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__I
timestamp 1669390400
transform -1 0 6608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__745__I
timestamp 1669390400
transform 1 0 63840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__I
timestamp 1669390400
transform 1 0 116480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__I
timestamp 1669390400
transform 1 0 75600 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__748__I
timestamp 1669390400
transform 1 0 81648 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__749__I
timestamp 1669390400
transform 1 0 46816 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__750__I
timestamp 1669390400
transform -1 0 116928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__I
timestamp 1669390400
transform 1 0 45584 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__752__I
timestamp 1669390400
transform 1 0 117824 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__753__I
timestamp 1669390400
transform -1 0 59808 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__754__I
timestamp 1669390400
transform -1 0 51968 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__755__I
timestamp 1669390400
transform 1 0 62608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__756__I
timestamp 1669390400
transform 1 0 79408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__757__I
timestamp 1669390400
transform 1 0 116480 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__758__I
timestamp 1669390400
transform 1 0 48720 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__759__I
timestamp 1669390400
transform 1 0 52192 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__760__I
timestamp 1669390400
transform 1 0 57680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__761__I
timestamp 1669390400
transform 1 0 40208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__762__I
timestamp 1669390400
transform -1 0 53760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__763__I
timestamp 1669390400
transform 1 0 71680 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__764__I
timestamp 1669390400
transform 1 0 71232 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__765__I
timestamp 1669390400
transform 1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__766__I
timestamp 1669390400
transform 1 0 49392 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__767__I
timestamp 1669390400
transform 1 0 88480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__768__I
timestamp 1669390400
transform 1 0 42896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__769__I
timestamp 1669390400
transform 1 0 71120 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__770__I
timestamp 1669390400
transform -1 0 68768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__771__I
timestamp 1669390400
transform 1 0 70112 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1669390400
transform -1 0 87920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 63168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 75040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 55216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 66864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 62160 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 65744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 67424 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1669390400
transform 1 0 82992 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout239_I
timestamp 1669390400
transform 1 0 12320 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout240_I
timestamp 1669390400
transform -1 0 22848 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout241_I
timestamp 1669390400
transform 1 0 114352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout242_I
timestamp 1669390400
transform -1 0 68208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout243_I
timestamp 1669390400
transform 1 0 62944 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 60032 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 117152 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 36960 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 49616 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform 1 0 116928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 41552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 57680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform 1 0 1680 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 114464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 1904 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 116816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 75712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform -1 0 56112 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform 1 0 17360 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 9968 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform 1 0 48720 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform 1 0 56560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform -1 0 1904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform -1 0 1904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform -1 0 1904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform 1 0 2128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1669390400
transform 1 0 117824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1669390400
transform -1 0 43792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1669390400
transform 1 0 116816 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1669390400
transform -1 0 21280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1669390400
transform 1 0 33040 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1669390400
transform -1 0 45136 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1669390400
transform -1 0 70448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1669390400
transform 1 0 116816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1669390400
transform 1 0 37408 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1669390400
transform -1 0 108752 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1669390400
transform 1 0 2352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1669390400
transform 1 0 5712 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1669390400
transform 1 0 63952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1669390400
transform -1 0 1904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1669390400
transform -1 0 1904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1669390400
transform -1 0 1904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1669390400
transform 1 0 45360 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1669390400
transform -1 0 1904 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1669390400
transform -1 0 53200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1669390400
transform -1 0 1904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1669390400
transform -1 0 95984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1669390400
transform -1 0 1904 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1669390400
transform -1 0 117152 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1669390400
transform -1 0 118048 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1669390400
transform -1 0 92624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1669390400
transform -1 0 40880 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1669390400
transform 1 0 117264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1669390400
transform -1 0 81200 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1669390400
transform -1 0 117152 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1669390400
transform -1 0 91392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1669390400
transform 1 0 106848 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1669390400
transform 1 0 116816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1669390400
transform -1 0 72240 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1669390400
transform -1 0 110992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1669390400
transform -1 0 1904 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1669390400
transform -1 0 14672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1669390400
transform 1 0 116816 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1669390400
transform -1 0 118048 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1669390400
transform -1 0 29456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1669390400
transform -1 0 114240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1669390400
transform -1 0 1904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1669390400
transform -1 0 22064 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1669390400
transform -1 0 38192 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1669390400
transform 1 0 116816 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1669390400
transform -1 0 1904 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1669390400
transform 1 0 2352 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1669390400
transform 1 0 1680 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1669390400
transform 1 0 5152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1669390400
transform 1 0 2128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1669390400
transform -1 0 117152 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1669390400
transform -1 0 69104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1669390400
transform -1 0 81872 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1669390400
transform -1 0 110992 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1669390400
transform -1 0 5936 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1669390400
transform -1 0 18032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1669390400
transform -1 0 1904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1669390400
transform -1 0 114912 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1669390400
transform -1 0 1904 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1669390400
transform -1 0 117152 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1669390400
transform -1 0 117152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1669390400
transform -1 0 83552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1669390400
transform -1 0 99232 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1669390400
transform -1 0 28784 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1669390400
transform -1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1669390400
transform -1 0 117152 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1669390400
transform -1 0 98000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1669390400
transform -1 0 117152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1669390400
transform -1 0 1904 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1669390400
transform -1 0 117152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1669390400
transform 1 0 21504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1669390400
transform -1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1669390400
transform 1 0 116816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1669390400
transform 1 0 95088 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1669390400
transform 1 0 116816 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1669390400
transform -1 0 116816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1669390400
transform 1 0 1680 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1669390400
transform -1 0 12880 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1669390400
transform -1 0 86576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1669390400
transform 1 0 1680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1669390400
transform -1 0 1904 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1669390400
transform -1 0 115920 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output142_I
timestamp 1669390400
transform 1 0 3472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output143_I
timestamp 1669390400
transform 1 0 114352 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output144_I
timestamp 1669390400
transform -1 0 114576 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output145_I
timestamp 1669390400
transform -1 0 117600 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1669390400
transform 1 0 3472 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1669390400
transform 1 0 49168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1669390400
transform -1 0 114576 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1669390400
transform 1 0 15344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1669390400
transform 1 0 100240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1669390400
transform 1 0 78288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1669390400
transform 1 0 9632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1669390400
transform 1 0 81648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1669390400
transform 1 0 57344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output155_I
timestamp 1669390400
transform -1 0 43344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output156_I
timestamp 1669390400
transform 1 0 3472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output157_I
timestamp 1669390400
transform 1 0 87920 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output158_I
timestamp 1669390400
transform 1 0 56448 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output159_I
timestamp 1669390400
transform 1 0 49392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output160_I
timestamp 1669390400
transform 1 0 85232 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output161_I
timestamp 1669390400
transform -1 0 88592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output162_I
timestamp 1669390400
transform -1 0 76496 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1669390400
transform 1 0 112336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output164_I
timestamp 1669390400
transform 1 0 110768 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1669390400
transform 1 0 114352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1669390400
transform 1 0 100464 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output167_I
timestamp 1669390400
transform 1 0 114352 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output168_I
timestamp 1669390400
transform 1 0 5600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output169_I
timestamp 1669390400
transform 1 0 3472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output170_I
timestamp 1669390400
transform -1 0 3696 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output171_I
timestamp 1669390400
transform 1 0 75488 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output172_I
timestamp 1669390400
transform 1 0 32816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output173_I
timestamp 1669390400
transform -1 0 3696 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output174_I
timestamp 1669390400
transform 1 0 35504 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output176_I
timestamp 1669390400
transform -1 0 3696 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output178_I
timestamp 1669390400
transform -1 0 59248 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output179_I
timestamp 1669390400
transform 1 0 52752 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output180_I
timestamp 1669390400
transform -1 0 63056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output181_I
timestamp 1669390400
transform -1 0 114576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output182_I
timestamp 1669390400
transform -1 0 116816 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output183_I
timestamp 1669390400
transform 1 0 3696 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output184_I
timestamp 1669390400
transform 1 0 114352 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output185_I
timestamp 1669390400
transform 1 0 36512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output186_I
timestamp 1669390400
transform -1 0 114576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output187_I
timestamp 1669390400
transform -1 0 3696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output188_I
timestamp 1669390400
transform -1 0 114576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output190_I
timestamp 1669390400
transform -1 0 114576 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output192_I
timestamp 1669390400
transform -1 0 3696 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output193_I
timestamp 1669390400
transform 1 0 114352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output194_I
timestamp 1669390400
transform 1 0 3472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output195_I
timestamp 1669390400
transform 1 0 71232 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output199_I
timestamp 1669390400
transform -1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output201_I
timestamp 1669390400
transform -1 0 114576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output203_I
timestamp 1669390400
transform -1 0 114576 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output204_I
timestamp 1669390400
transform -1 0 114128 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output205_I
timestamp 1669390400
transform 1 0 46928 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1669390400
transform 1 0 114352 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1669390400
transform 1 0 3472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output208_I
timestamp 1669390400
transform 1 0 114352 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output209_I
timestamp 1669390400
transform 1 0 6048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output210_I
timestamp 1669390400
transform 1 0 116592 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output211_I
timestamp 1669390400
transform 1 0 91168 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1669390400
transform -1 0 114576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output213_I
timestamp 1669390400
transform -1 0 85904 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output214_I
timestamp 1669390400
transform -1 0 3696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output215_I
timestamp 1669390400
transform 1 0 3472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output216_I
timestamp 1669390400
transform 1 0 80528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output217_I
timestamp 1669390400
transform -1 0 3696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1669390400
transform -1 0 94864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output219_I
timestamp 1669390400
transform 1 0 3472 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output220_I
timestamp 1669390400
transform -1 0 3696 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output221_I
timestamp 1669390400
transform -1 0 33712 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output222_I
timestamp 1669390400
transform -1 0 3696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output223_I
timestamp 1669390400
transform -1 0 26992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output224_I
timestamp 1669390400
transform 1 0 10528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output225_I
timestamp 1669390400
transform 1 0 64400 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output226_I
timestamp 1669390400
transform 1 0 36624 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output227_I
timestamp 1669390400
transform 1 0 65296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output228_I
timestamp 1669390400
transform 1 0 84112 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output230_I
timestamp 1669390400
transform 1 0 3472 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output231_I
timestamp 1669390400
transform 1 0 114352 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output232_I
timestamp 1669390400
transform 1 0 28112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output233_I
timestamp 1669390400
transform -1 0 46256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output234_I
timestamp 1669390400
transform 1 0 3472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output235_I
timestamp 1669390400
transform 1 0 116928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1669390400
transform -1 0 73248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1669390400
transform 1 0 80528 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1669390400
transform 1 0 77840 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7
timestamp 1669390400
transform 1 0 2128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15
timestamp 1669390400
transform 1 0 3024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17
timestamp 1669390400
transform 1 0 3248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52
timestamp 1669390400
transform 1 0 7168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54
timestamp 1669390400
transform 1 0 7392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87
timestamp 1669390400
transform 1 0 11088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89
timestamp 1669390400
transform 1 0 11312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115
timestamp 1669390400
transform 1 0 14224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119
timestamp 1669390400
transform 1 0 14672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137
timestamp 1669390400
transform 1 0 16688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_194
timestamp 1669390400
transform 1 0 23072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_202 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_206
timestamp 1669390400
transform 1 0 24416 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_229
timestamp 1669390400
transform 1 0 26992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_233
timestamp 1669390400
transform 1 0 27440 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_238
timestamp 1669390400
transform 1 0 28000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_251
timestamp 1669390400
transform 1 0 29456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_269
timestamp 1669390400
transform 1 0 31472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_277
timestamp 1669390400
transform 1 0 32368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_287
timestamp 1669390400
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_295
timestamp 1669390400
transform 1 0 34384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_299
timestamp 1669390400
transform 1 0 34832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_323
timestamp 1669390400
transform 1 0 37520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_341
timestamp 1669390400
transform 1 0 39536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_356
timestamp 1669390400
transform 1 0 41216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1669390400
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_377
timestamp 1669390400
transform 1 0 43568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_407
timestamp 1669390400
transform 1 0 46928 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_415
timestamp 1669390400
transform 1 0 47824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_437
timestamp 1669390400
transform 1 0 50288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_463
timestamp 1669390400
transform 1 0 53200 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_471
timestamp 1669390400
transform 1 0 54096 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_495
timestamp 1669390400
transform 1 0 56784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_499
timestamp 1669390400
transform 1 0 57232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_503
timestamp 1669390400
transform 1 0 57680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_521
timestamp 1669390400
transform 1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_564
timestamp 1669390400
transform 1 0 64512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_579
timestamp 1669390400
transform 1 0 66192 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_601
timestamp 1669390400
transform 1 0 68656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_605
timestamp 1669390400
transform 1 0 69104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_623
timestamp 1669390400
transform 1 0 71120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_627
timestamp 1669390400
transform 1 0 71568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1669390400
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_642
timestamp 1669390400
transform 1 0 73248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_646
timestamp 1669390400
transform 1 0 73696 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_672
timestamp 1669390400
transform 1 0 76608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_676
timestamp 1669390400
transform 1 0 77056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_678
timestamp 1669390400
transform 1 0 77280 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_693
timestamp 1669390400
transform 1 0 78960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_697
timestamp 1669390400
transform 1 0 79408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_699
timestamp 1669390400
transform 1 0 79632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1669390400
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_707
timestamp 1669390400
transform 1 0 80528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_723
timestamp 1669390400
transform 1 0 82320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_731
timestamp 1669390400
transform 1 0 83216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_734
timestamp 1669390400
transform 1 0 83552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_737
timestamp 1669390400
transform 1 0 83888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_754
timestamp 1669390400
transform 1 0 85792 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_772
timestamp 1669390400
transform 1 0 87808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_776
timestamp 1669390400
transform 1 0 88256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_779
timestamp 1669390400
transform 1 0 88592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_795
timestamp 1669390400
transform 1 0 90384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_799
timestamp 1669390400
transform 1 0 90832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_801
timestamp 1669390400
transform 1 0 91056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_804
timestamp 1669390400
transform 1 0 91392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1669390400
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_824
timestamp 1669390400
transform 1 0 93632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_832
timestamp 1669390400
transform 1 0 94528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_835
timestamp 1669390400
transform 1 0 94864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1669390400
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_842
timestamp 1669390400
transform 1 0 95648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_845
timestamp 1669390400
transform 1 0 95984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_863
timestamp 1669390400
transform 1 0 98000 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_871
timestamp 1669390400
transform 1 0 98896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1669390400
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_892
timestamp 1669390400
transform 1 0 101248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_908
timestamp 1669390400
transform 1 0 103040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1669390400
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_927
timestamp 1669390400
transform 1 0 105168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_933
timestamp 1669390400
transform 1 0 105840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_941
timestamp 1669390400
transform 1 0 106736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_947
timestamp 1669390400
transform 1 0 107408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_955
timestamp 1669390400
transform 1 0 108304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_959
timestamp 1669390400
transform 1 0 108752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_965
timestamp 1669390400
transform 1 0 109424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_971
timestamp 1669390400
transform 1 0 110096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_975
timestamp 1669390400
transform 1 0 110544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1669390400
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1669390400
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_999
timestamp 1669390400
transform 1 0 113232 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1003
timestamp 1669390400
transform 1 0 113680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1005
timestamp 1669390400
transform 1 0 113904 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1008
timestamp 1669390400
transform 1 0 114240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1012
timestamp 1669390400
transform 1 0 114688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1669390400
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1669390400
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1034
timestamp 1669390400
transform 1 0 117152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1038
timestamp 1669390400
transform 1 0 117600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1044
timestamp 1669390400
transform 1 0 118272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_19
timestamp 1669390400
transform 1 0 3472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_35
timestamp 1669390400
transform 1 0 5264 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_43
timestamp 1669390400
transform 1 0 6160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_47
timestamp 1669390400
transform 1 0 6608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_63
timestamp 1669390400
transform 1 0 8400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_67
timestamp 1669390400
transform 1 0 8848 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_76
timestamp 1669390400
transform 1 0 9856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_80
timestamp 1669390400
transform 1 0 10304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1669390400
transform 1 0 10752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_92
timestamp 1669390400
transform 1 0 11648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_96
timestamp 1669390400
transform 1 0 12096 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_104
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_108
timestamp 1669390400
transform 1 0 13440 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_123
timestamp 1669390400
transform 1 0 15120 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_127
timestamp 1669390400
transform 1 0 15568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1669390400
transform 1 0 16464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_139
timestamp 1669390400
transform 1 0 16912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_146
timestamp 1669390400
transform 1 0 17696 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_149
timestamp 1669390400
transform 1 0 18032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_167
timestamp 1669390400
transform 1 0 20048 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_175
timestamp 1669390400
transform 1 0 20944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_178
timestamp 1669390400
transform 1 0 21280 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_182
timestamp 1669390400
transform 1 0 21728 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_198
timestamp 1669390400
transform 1 0 23520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1669390400
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_210
timestamp 1669390400
transform 1 0 24864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_237
timestamp 1669390400
transform 1 0 27888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_241
timestamp 1669390400
transform 1 0 28336 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_257
timestamp 1669390400
transform 1 0 30128 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_302
timestamp 1669390400
transform 1 0 35168 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_310
timestamp 1669390400
transform 1 0 36064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_316
timestamp 1669390400
transform 1 0 36736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_320
timestamp 1669390400
transform 1 0 37184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_322
timestamp 1669390400
transform 1 0 37408 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_325
timestamp 1669390400
transform 1 0 37744 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_341
timestamp 1669390400
transform 1 0 39536 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_349
timestamp 1669390400
transform 1 0 40432 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_353
timestamp 1669390400
transform 1 0 40880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_361
timestamp 1669390400
transform 1 0 41776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_377
timestamp 1669390400
transform 1 0 43568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_395
timestamp 1669390400
transform 1 0 45584 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_403
timestamp 1669390400
transform 1 0 46480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_407
timestamp 1669390400
transform 1 0 46928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_423
timestamp 1669390400
transform 1 0 48720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_431
timestamp 1669390400
transform 1 0 49616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_437
timestamp 1669390400
transform 1 0 50288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_445
timestamp 1669390400
transform 1 0 51184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_461
timestamp 1669390400
transform 1 0 52976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_479
timestamp 1669390400
transform 1 0 54992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1669390400
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_502
timestamp 1669390400
transform 1 0 57568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_506
timestamp 1669390400
transform 1 0 58016 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_521
timestamp 1669390400
transform 1 0 59696 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_539
timestamp 1669390400
transform 1 0 61712 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_547
timestamp 1669390400
transform 1 0 62608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_551
timestamp 1669390400
transform 1 0 63056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1669390400
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_573
timestamp 1669390400
transform 1 0 65520 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_589
timestamp 1669390400
transform 1 0 67312 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_591
timestamp 1669390400
transform 1 0 67536 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_598
timestamp 1669390400
transform 1 0 68320 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_602
timestamp 1669390400
transform 1 0 68768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_610
timestamp 1669390400
transform 1 0 69664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_614
timestamp 1669390400
transform 1 0 70112 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_617
timestamp 1669390400
transform 1 0 70448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_635
timestamp 1669390400
transform 1 0 72464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_656
timestamp 1669390400
transform 1 0 74816 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_666
timestamp 1669390400
transform 1 0 75936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_672
timestamp 1669390400
transform 1 0 76608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_680
timestamp 1669390400
transform 1 0 77504 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_684
timestamp 1669390400
transform 1 0 77952 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_686
timestamp 1669390400
transform 1 0 78176 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_689
timestamp 1669390400
transform 1 0 78512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_705
timestamp 1669390400
transform 1 0 80304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1669390400
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_712
timestamp 1669390400
transform 1 0 81088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_716
timestamp 1669390400
transform 1 0 81536 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_719
timestamp 1669390400
transform 1 0 81872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_735
timestamp 1669390400
transform 1 0 83664 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_751
timestamp 1669390400
transform 1 0 85456 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_761
timestamp 1669390400
transform 1 0 86576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_779
timestamp 1669390400
transform 1 0 88592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_783
timestamp 1669390400
transform 1 0 89040 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_799
timestamp 1669390400
transform 1 0 90832 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_807
timestamp 1669390400
transform 1 0 91728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_811
timestamp 1669390400
transform 1 0 92176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_815
timestamp 1669390400
transform 1 0 92624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_833
timestamp 1669390400
transform 1 0 94640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_849
timestamp 1669390400
transform 1 0 96432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1669390400
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_854
timestamp 1669390400
transform 1 0 96992 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_858
timestamp 1669390400
transform 1 0 97440 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_860
timestamp 1669390400
transform 1 0 97664 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_863
timestamp 1669390400
transform 1 0 98000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_881
timestamp 1669390400
transform 1 0 100016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_885
timestamp 1669390400
transform 1 0 100464 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_893
timestamp 1669390400
transform 1 0 101360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_909
timestamp 1669390400
transform 1 0 103152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_917
timestamp 1669390400
transform 1 0 104048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_921
timestamp 1669390400
transform 1 0 104496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_925 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 104944 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_957
timestamp 1669390400
transform 1 0 108528 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_973
timestamp 1669390400
transform 1 0 110320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_977
timestamp 1669390400
transform 1 0 110768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1669390400
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1669390400
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1011
timestamp 1669390400
transform 1 0 114576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1029
timestamp 1669390400
transform 1 0 116592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1031
timestamp 1669390400
transform 1 0 116816 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1038
timestamp 1669390400
transform 1 0 117600 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1042
timestamp 1669390400
transform 1 0 118048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1044
timestamp 1669390400
transform 1 0 118272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_17
timestamp 1669390400
transform 1 0 3248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1669390400
transform 1 0 5040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_40
timestamp 1669390400
transform 1 0 5824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_44
timestamp 1669390400
transform 1 0 6272 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_76
timestamp 1669390400
transform 1 0 9856 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_92
timestamp 1669390400
transform 1 0 11648 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_100
timestamp 1669390400
transform 1 0 12544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_104
timestamp 1669390400
transform 1 0 12992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_225
timestamp 1669390400
transform 1 0 26544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_229
timestamp 1669390400
transform 1 0 26992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_245
timestamp 1669390400
transform 1 0 28784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_337
timestamp 1669390400
transform 1 0 39088 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_345
timestamp 1669390400
transform 1 0 39984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_363
timestamp 1669390400
transform 1 0 42000 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_371
timestamp 1669390400
transform 1 0 42896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_375
timestamp 1669390400
transform 1 0 43344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_379
timestamp 1669390400
transform 1 0 43792 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_387
timestamp 1669390400
transform 1 0 44688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_396
timestamp 1669390400
transform 1 0 45696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_398
timestamp 1669390400
transform 1 0 45920 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_401
timestamp 1669390400
transform 1 0 46256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_417
timestamp 1669390400
transform 1 0 48048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_425
timestamp 1669390400
transform 1 0 48944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_429
timestamp 1669390400
transform 1 0 49392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_439
timestamp 1669390400
transform 1 0 50512 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_455
timestamp 1669390400
transform 1 0 52304 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_459
timestamp 1669390400
transform 1 0 52752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_471
timestamp 1669390400
transform 1 0 54096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_479
timestamp 1669390400
transform 1 0 54992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_483
timestamp 1669390400
transform 1 0 55440 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_515
timestamp 1669390400
transform 1 0 59024 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_519
timestamp 1669390400
transform 1 0 59472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_523
timestamp 1669390400
transform 1 0 59920 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1669390400
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_550
timestamp 1669390400
transform 1 0 62944 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_558
timestamp 1669390400
transform 1 0 63840 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_561
timestamp 1669390400
transform 1 0 64176 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_593
timestamp 1669390400
transform 1 0 67760 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_601
timestamp 1669390400
transform 1 0 68656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_669
timestamp 1669390400
transform 1 0 76272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1669390400
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_740
timestamp 1669390400
transform 1 0 84224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1669390400
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_747
timestamp 1669390400
transform 1 0 85008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_811
timestamp 1669390400
transform 1 0 92176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1669390400
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_818
timestamp 1669390400
transform 1 0 92960 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_850
timestamp 1669390400
transform 1 0 96544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_866
timestamp 1669390400
transform 1 0 98336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_870
timestamp 1669390400
transform 1 0 98784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_878
timestamp 1669390400
transform 1 0 99680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_882
timestamp 1669390400
transform 1 0 100128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1669390400
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_889
timestamp 1669390400
transform 1 0 100912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_895
timestamp 1669390400
transform 1 0 101584 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_927
timestamp 1669390400
transform 1 0 105168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_943
timestamp 1669390400
transform 1 0 106960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_951
timestamp 1669390400
transform 1 0 107856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_955
timestamp 1669390400
transform 1 0 108304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1669390400
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_960
timestamp 1669390400
transform 1 0 108864 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_976
timestamp 1669390400
transform 1 0 110656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_980
timestamp 1669390400
transform 1 0 111104 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_984
timestamp 1669390400
transform 1 0 111552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_992
timestamp 1669390400
transform 1 0 112448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1010
timestamp 1669390400
transform 1 0 114464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1669390400
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1669390400
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1034
timestamp 1669390400
transform 1 0 117152 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1042
timestamp 1669390400
transform 1 0 118048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1044
timestamp 1669390400
transform 1 0 118272 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_17
timestamp 1669390400
transform 1 0 3248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_21
timestamp 1669390400
transform 1 0 3696 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_29
timestamp 1669390400
transform 1 0 4592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_33
timestamp 1669390400
transform 1 0 5040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_36
timestamp 1669390400
transform 1 0 5376 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_68
timestamp 1669390400
transform 1 0 8960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_361
timestamp 1669390400
transform 1 0 41776 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_365
timestamp 1669390400
transform 1 0 42224 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_397
timestamp 1669390400
transform 1 0 45808 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1669390400
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_419
timestamp 1669390400
transform 1 0 48272 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_423
timestamp 1669390400
transform 1 0 48720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_705
timestamp 1669390400
transform 1 0 80304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1669390400
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_712
timestamp 1669390400
transform 1 0 81088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_776
timestamp 1669390400
transform 1 0 88256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1669390400
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1669390400
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_847
timestamp 1669390400
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1669390400
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_854
timestamp 1669390400
transform 1 0 96992 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_918
timestamp 1669390400
transform 1 0 104160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1669390400
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_925
timestamp 1669390400
transform 1 0 104944 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_989
timestamp 1669390400
transform 1 0 112112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1669390400
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_996
timestamp 1669390400
transform 1 0 112896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1011
timestamp 1669390400
transform 1 0 114576 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1029
timestamp 1669390400
transform 1 0 116592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1033
timestamp 1669390400
transform 1 0 117040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1037
timestamp 1669390400
transform 1 0 117488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_17
timestamp 1669390400
transform 1 0 3248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_21
timestamp 1669390400
transform 1 0 3696 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_29
timestamp 1669390400
transform 1 0 4592 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_33
timestamp 1669390400
transform 1 0 5040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1669390400
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1669390400
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1669390400
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1669390400
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1669390400
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1669390400
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_818
timestamp 1669390400
transform 1 0 92960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_882
timestamp 1669390400
transform 1 0 100128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1669390400
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_889
timestamp 1669390400
transform 1 0 100912 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1669390400
transform 1 0 108080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1669390400
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_960
timestamp 1669390400
transform 1 0 108864 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_992
timestamp 1669390400
transform 1 0 112448 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1008
timestamp 1669390400
transform 1 0 114240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1028
timestamp 1669390400
transform 1 0 116480 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1031
timestamp 1669390400
transform 1 0 116816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1038
timestamp 1669390400
transform 1 0 117600 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1042
timestamp 1669390400
transform 1 0 118048 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1044
timestamp 1669390400
transform 1 0 118272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_7
timestamp 1669390400
transform 1 0 2128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_11
timestamp 1669390400
transform 1 0 2576 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_43
timestamp 1669390400
transform 1 0 6160 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_59
timestamp 1669390400
transform 1 0 7952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_67
timestamp 1669390400
transform 1 0 8848 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1669390400
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1669390400
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1669390400
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1669390400
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1669390400
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1669390400
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1669390400
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1669390400
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_854
timestamp 1669390400
transform 1 0 96992 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_918
timestamp 1669390400
transform 1 0 104160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1669390400
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1669390400
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1669390400
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1669390400
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_996
timestamp 1669390400
transform 1 0 112896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1012
timestamp 1669390400
transform 1 0 114688 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1027
timestamp 1669390400
transform 1 0 116368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1031
timestamp 1669390400
transform 1 0 116816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1039
timestamp 1669390400
transform 1 0 117712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1043
timestamp 1669390400
transform 1 0 118160 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_550
timestamp 1669390400
transform 1 0 62944 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_560
timestamp 1669390400
transform 1 0 64064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_568
timestamp 1669390400
transform 1 0 64960 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_600
timestamp 1669390400
transform 1 0 68544 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1669390400
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1669390400
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1669390400
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1669390400
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1669390400
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1669390400
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1669390400
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1669390400
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1669390400
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1669390400
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1669390400
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_960
timestamp 1669390400
transform 1 0 108864 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_992
timestamp 1669390400
transform 1 0 112448 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1008
timestamp 1669390400
transform 1 0 114240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1011
timestamp 1669390400
transform 1 0 114576 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1027
timestamp 1669390400
transform 1 0 116368 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1031
timestamp 1669390400
transform 1 0 116816 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1039
timestamp 1669390400
transform 1 0 117712 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1043
timestamp 1669390400
transform 1 0 118160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1669390400
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1669390400
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1669390400
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1669390400
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1669390400
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1669390400
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1669390400
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1669390400
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1669390400
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1669390400
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1669390400
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1669390400
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1669390400
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1669390400
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_996
timestamp 1669390400
transform 1 0 112896 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1028
timestamp 1669390400
transform 1 0 116480 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_1032
timestamp 1669390400
transform 1 0 116928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1040
timestamp 1669390400
transform 1 0 117824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1044
timestamp 1669390400
transform 1 0 118272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1669390400
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1669390400
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1669390400
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1669390400
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1669390400
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1669390400
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1669390400
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1669390400
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1669390400
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1669390400
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1669390400
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_960
timestamp 1669390400
transform 1 0 108864 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_992
timestamp 1669390400
transform 1 0 112448 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1008
timestamp 1669390400
transform 1 0 114240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1012
timestamp 1669390400
transform 1 0 114688 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1027
timestamp 1669390400
transform 1 0 116368 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1031
timestamp 1669390400
transform 1 0 116816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1038
timestamp 1669390400
transform 1 0 117600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1042
timestamp 1669390400
transform 1 0 118048 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1044
timestamp 1669390400
transform 1 0 118272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_17
timestamp 1669390400
transform 1 0 3248 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_21
timestamp 1669390400
transform 1 0 3696 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_53
timestamp 1669390400
transform 1 0 7280 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1669390400
transform 1 0 9072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1669390400
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1669390400
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1669390400
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1669390400
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1669390400
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1669390400
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1669390400
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1669390400
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1669390400
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1669390400
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1669390400
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1669390400
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1669390400
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1669390400
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_996
timestamp 1669390400
transform 1 0 112896 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1028
timestamp 1669390400
transform 1 0 116480 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1044
timestamp 1669390400
transform 1 0 118272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_6
timestamp 1669390400
transform 1 0 2016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_8
timestamp 1669390400
transform 1 0 2240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_15
timestamp 1669390400
transform 1 0 3024 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_19
timestamp 1669390400
transform 1 0 3472 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1669390400
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1669390400
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1669390400
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1669390400
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1669390400
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1669390400
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1669390400
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1669390400
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1669390400
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1669390400
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1669390400
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1669390400
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1669390400
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1669390400
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_1031
timestamp 1669390400
transform 1 0 116816 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1039
timestamp 1669390400
transform 1 0 117712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1043
timestamp 1669390400
transform 1 0 118160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_17
timestamp 1669390400
transform 1 0 3248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_49
timestamp 1669390400
transform 1 0 6832 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_65
timestamp 1669390400
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1669390400
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1669390400
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1669390400
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1669390400
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1669390400
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1669390400
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1669390400
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1669390400
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1669390400
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1669390400
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1669390400
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1669390400
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1669390400
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1669390400
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1669390400
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_996
timestamp 1669390400
transform 1 0 112896 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1012
timestamp 1669390400
transform 1 0 114688 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_1029
timestamp 1669390400
transform 1 0 116592 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_1033
timestamp 1669390400
transform 1 0 117040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1041
timestamp 1669390400
transform 1 0 117936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1669390400
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1669390400
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1669390400
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1669390400
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1669390400
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1669390400
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1669390400
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1669390400
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1669390400
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1669390400
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1669390400
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1669390400
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1669390400
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1669390400
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_1031
timestamp 1669390400
transform 1 0 116816 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1039
timestamp 1669390400
transform 1 0 117712 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1043
timestamp 1669390400
transform 1 0 118160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1669390400
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1669390400
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1669390400
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1669390400
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1669390400
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1669390400
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1669390400
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1669390400
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1669390400
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1669390400
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1669390400
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1669390400
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1669390400
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1669390400
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_996
timestamp 1669390400
transform 1 0 112896 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_1028
timestamp 1669390400
transform 1 0 116480 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1044
timestamp 1669390400
transform 1 0 118272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1669390400
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1669390400
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1669390400
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1669390400
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1669390400
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1669390400
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1669390400
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1669390400
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1669390400
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1669390400
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1669390400
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_960
timestamp 1669390400
transform 1 0 108864 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_992
timestamp 1669390400
transform 1 0 112448 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1008
timestamp 1669390400
transform 1 0 114240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1011
timestamp 1669390400
transform 1 0 114576 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1027
timestamp 1669390400
transform 1 0 116368 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_1031
timestamp 1669390400
transform 1 0 116816 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1039
timestamp 1669390400
transform 1 0 117712 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1043
timestamp 1669390400
transform 1 0 118160 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_460
timestamp 1669390400
transform 1 0 52864 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_464
timestamp 1669390400
transform 1 0 53312 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_468
timestamp 1669390400
transform 1 0 53760 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_476
timestamp 1669390400
transform 1 0 54656 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1669390400
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1669390400
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1669390400
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1669390400
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1669390400
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1669390400
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1669390400
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1669390400
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1669390400
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1669390400
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1669390400
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1669390400
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1669390400
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1669390400
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_996
timestamp 1669390400
transform 1 0 112896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1004
timestamp 1669390400
transform 1 0 113792 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1008
timestamp 1669390400
transform 1 0 114240 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1011
timestamp 1669390400
transform 1 0 114576 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_1027
timestamp 1669390400
transform 1 0 116368 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1043
timestamp 1669390400
transform 1 0 118160 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1669390400
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1669390400
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1669390400
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1669390400
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1669390400
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1669390400
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1669390400
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1669390400
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1669390400
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1669390400
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1669390400
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1669390400
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1669390400
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1669390400
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1031
timestamp 1669390400
transform 1 0 116816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1039
timestamp 1669390400
transform 1 0 117712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1043
timestamp 1669390400
transform 1 0 118160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_17
timestamp 1669390400
transform 1 0 3248 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_21
timestamp 1669390400
transform 1 0 3696 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_53
timestamp 1669390400
transform 1 0 7280 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_69
timestamp 1669390400
transform 1 0 9072 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1669390400
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1669390400
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1669390400
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1669390400
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1669390400
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1669390400
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1669390400
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1669390400
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1669390400
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1669390400
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1669390400
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1669390400
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1669390400
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1669390400
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_996
timestamp 1669390400
transform 1 0 112896 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_1028
timestamp 1669390400
transform 1 0 116480 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1036
timestamp 1669390400
transform 1 0 117376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1044
timestamp 1669390400
transform 1 0 118272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_7
timestamp 1669390400
transform 1 0 2128 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_23
timestamp 1669390400
transform 1 0 3920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_31
timestamp 1669390400
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1669390400
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1669390400
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1669390400
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1669390400
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1669390400
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1669390400
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1669390400
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1669390400
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1669390400
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1669390400
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1669390400
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1669390400
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1669390400
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1669390400
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_1031
timestamp 1669390400
transform 1 0 116816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1039
timestamp 1669390400
transform 1 0 117712 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_1043
timestamp 1669390400
transform 1 0 118160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_7
timestamp 1669390400
transform 1 0 2128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1669390400
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1669390400
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1669390400
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1669390400
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1669390400
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1669390400
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1669390400
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1669390400
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1669390400
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1669390400
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1669390400
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1669390400
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1669390400
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1669390400
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_996
timestamp 1669390400
transform 1 0 112896 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1028
timestamp 1669390400
transform 1 0 116480 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_1032
timestamp 1669390400
transform 1 0 116928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1040
timestamp 1669390400
transform 1 0 117824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1044
timestamp 1669390400
transform 1 0 118272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1669390400
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1669390400
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1669390400
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1669390400
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1669390400
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1669390400
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1669390400
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1669390400
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1669390400
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1669390400
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1669390400
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_960
timestamp 1669390400
transform 1 0 108864 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_992
timestamp 1669390400
transform 1 0 112448 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1008
timestamp 1669390400
transform 1 0 114240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1012
timestamp 1669390400
transform 1 0 114688 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1027
timestamp 1669390400
transform 1 0 116368 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1031
timestamp 1669390400
transform 1 0 116816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1038
timestamp 1669390400
transform 1 0 117600 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1042
timestamp 1669390400
transform 1 0 118048 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1044
timestamp 1669390400
transform 1 0 118272 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_389
timestamp 1669390400
transform 1 0 44912 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_395
timestamp 1669390400
transform 1 0 45584 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_412
timestamp 1669390400
transform 1 0 47488 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_416
timestamp 1669390400
transform 1 0 47936 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_420
timestamp 1669390400
transform 1 0 48384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_424
timestamp 1669390400
transform 1 0 48832 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1669390400
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1669390400
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1669390400
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1669390400
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1669390400
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1669390400
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1669390400
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1669390400
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1669390400
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1669390400
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1669390400
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1669390400
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1669390400
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1669390400
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_996
timestamp 1669390400
transform 1 0 112896 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_1028
timestamp 1669390400
transform 1 0 116480 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1044
timestamp 1669390400
transform 1 0 118272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_5
timestamp 1669390400
transform 1 0 1904 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_21
timestamp 1669390400
transform 1 0 3696 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_29
timestamp 1669390400
transform 1 0 4592 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_33
timestamp 1669390400
transform 1 0 5040 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_337
timestamp 1669390400
transform 1 0 39088 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_345
timestamp 1669390400
transform 1 0 39984 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_349
timestamp 1669390400
transform 1 0 40432 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_381
timestamp 1669390400
transform 1 0 44016 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_422
timestamp 1669390400
transform 1 0 48608 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_426
timestamp 1669390400
transform 1 0 49056 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_458
timestamp 1669390400
transform 1 0 52640 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1669390400
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1669390400
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_747
timestamp 1669390400
transform 1 0 85008 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_779
timestamp 1669390400
transform 1 0 88592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_787
timestamp 1669390400
transform 1 0 89488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_791
timestamp 1669390400
transform 1 0 89936 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_794
timestamp 1669390400
transform 1 0 90272 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_798
timestamp 1669390400
transform 1 0 90720 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1669390400
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_818
timestamp 1669390400
transform 1 0 92960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_821
timestamp 1669390400
transform 1 0 93296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_885
timestamp 1669390400
transform 1 0 100464 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1669390400
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1669390400
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1669390400
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1669390400
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1669390400
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1669390400
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_1031
timestamp 1669390400
transform 1 0 116816 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1039
timestamp 1669390400
transform 1 0 117712 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_1043
timestamp 1669390400
transform 1 0 118160 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_17
timestamp 1669390400
transform 1 0 3248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_21
timestamp 1669390400
transform 1 0 3696 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_53
timestamp 1669390400
transform 1 0 7280 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_69
timestamp 1669390400
transform 1 0 9072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_373
timestamp 1669390400
transform 1 0 43120 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_387
timestamp 1669390400
transform 1 0 44688 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_418
timestamp 1669390400
transform 1 0 48160 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_422
timestamp 1669390400
transform 1 0 48608 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1669390400
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1669390400
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1669390400
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1669390400
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1669390400
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_783
timestamp 1669390400
transform 1 0 89040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_791
timestamp 1669390400
transform 1 0 89936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_795
timestamp 1669390400
transform 1 0 90384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_799
timestamp 1669390400
transform 1 0 90832 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_830
timestamp 1669390400
transform 1 0 94304 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_846
timestamp 1669390400
transform 1 0 96096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_850
timestamp 1669390400
transform 1 0 96544 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1669390400
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1669390400
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1669390400
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1669390400
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1669390400
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1669390400
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_996
timestamp 1669390400
transform 1 0 112896 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_1028
timestamp 1669390400
transform 1 0 116480 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1044
timestamp 1669390400
transform 1 0 118272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_28
timestamp 1669390400
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_32
timestamp 1669390400
transform 1 0 4928 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_395
timestamp 1669390400
transform 1 0 45584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_412
timestamp 1669390400
transform 1 0 47488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_416
timestamp 1669390400
transform 1 0 47936 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_420
timestamp 1669390400
transform 1 0 48384 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_452
timestamp 1669390400
transform 1 0 51968 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_678
timestamp 1669390400
transform 1 0 77280 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_708
timestamp 1669390400
transform 1 0 80640 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1669390400
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1669390400
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_747
timestamp 1669390400
transform 1 0 85008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_779
timestamp 1669390400
transform 1 0 88592 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_795
timestamp 1669390400
transform 1 0 90384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_803
timestamp 1669390400
transform 1 0 91280 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_805
timestamp 1669390400
transform 1 0 91504 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_812
timestamp 1669390400
transform 1 0 92288 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1669390400
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1669390400
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1669390400
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1669390400
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1669390400
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1669390400
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_960
timestamp 1669390400
transform 1 0 108864 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_992
timestamp 1669390400
transform 1 0 112448 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1008
timestamp 1669390400
transform 1 0 114240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1012
timestamp 1669390400
transform 1 0 114688 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1027
timestamp 1669390400
transform 1 0 116368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_1031
timestamp 1669390400
transform 1 0 116816 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1039
timestamp 1669390400
transform 1 0 117712 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1043
timestamp 1669390400
transform 1 0 118160 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1669390400
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_21
timestamp 1669390400
transform 1 0 3696 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_53
timestamp 1669390400
transform 1 0 7280 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_69
timestamp 1669390400
transform 1 0 9072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_389
timestamp 1669390400
transform 1 0 44912 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_399
timestamp 1669390400
transform 1 0 46032 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_415
timestamp 1669390400
transform 1 0 47824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_423
timestamp 1669390400
transform 1 0 48720 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_673
timestamp 1669390400
transform 1 0 76720 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_677
timestamp 1669390400
transform 1 0 77168 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_685
timestamp 1669390400
transform 1 0 78064 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_702
timestamp 1669390400
transform 1 0 79968 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_706
timestamp 1669390400
transform 1 0 80416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1669390400
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1669390400
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1669390400
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1669390400
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1669390400
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1669390400
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1669390400
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1669390400
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1669390400
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1669390400
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1669390400
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1669390400
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_996
timestamp 1669390400
transform 1 0 112896 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1030
timestamp 1669390400
transform 1 0 116704 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1038
timestamp 1669390400
transform 1 0 117600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1042
timestamp 1669390400
transform 1 0 118048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1044
timestamp 1669390400
transform 1 0 118272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_409
timestamp 1669390400
transform 1 0 47152 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_413
timestamp 1669390400
transform 1 0 47600 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_417
timestamp 1669390400
transform 1 0 48048 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_449
timestamp 1669390400
transform 1 0 51632 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_457
timestamp 1669390400
transform 1 0 52528 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_680
timestamp 1669390400
transform 1 0 77504 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_682
timestamp 1669390400
transform 1 0 77728 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_685
timestamp 1669390400
transform 1 0 78064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_689
timestamp 1669390400
transform 1 0 78512 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_721
timestamp 1669390400
transform 1 0 82096 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_737
timestamp 1669390400
transform 1 0 83888 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1669390400
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1669390400
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1669390400
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1669390400
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1669390400
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1669390400
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1669390400
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1669390400
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1669390400
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1669390400
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1669390400
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1669390400
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_1031
timestamp 1669390400
transform 1 0 116816 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1039
timestamp 1669390400
transform 1 0 117712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1043
timestamp 1669390400
transform 1 0 118160 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_17
timestamp 1669390400
transform 1 0 3248 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_21
timestamp 1669390400
transform 1 0 3696 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_53
timestamp 1669390400
transform 1 0 7280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_69
timestamp 1669390400
transform 1 0 9072 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_373
timestamp 1669390400
transform 1 0 43120 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_381
timestamp 1669390400
transform 1 0 44016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_385
timestamp 1669390400
transform 1 0 44464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_415
timestamp 1669390400
transform 1 0 47824 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_419
timestamp 1669390400
transform 1 0 48272 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_423
timestamp 1669390400
transform 1 0 48720 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1669390400
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1669390400
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1669390400
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1669390400
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1669390400
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1669390400
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1669390400
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1669390400
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1669390400
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1669390400
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1669390400
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1669390400
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1669390400
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1669390400
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_996
timestamp 1669390400
transform 1 0 112896 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_1028
timestamp 1669390400
transform 1 0 116480 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1044
timestamp 1669390400
transform 1 0 118272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_19
timestamp 1669390400
transform 1 0 3472 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_399
timestamp 1669390400
transform 1 0 46032 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_431
timestamp 1669390400
transform 1 0 49616 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_447
timestamp 1669390400
transform 1 0 51408 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_455
timestamp 1669390400
transform 1 0 52304 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_459
timestamp 1669390400
transform 1 0 52752 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1669390400
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1669390400
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1669390400
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1669390400
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1669390400
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1669390400
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1669390400
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1669390400
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1669390400
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1669390400
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1669390400
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1669390400
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1669390400
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1669390400
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_1031
timestamp 1669390400
transform 1 0 116816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1039
timestamp 1669390400
transform 1 0 117712 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_1043
timestamp 1669390400
transform 1 0 118160 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_5
timestamp 1669390400
transform 1 0 1904 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_9
timestamp 1669390400
transform 1 0 2352 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_41
timestamp 1669390400
transform 1 0 5936 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_57
timestamp 1669390400
transform 1 0 7728 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_65
timestamp 1669390400
transform 1 0 8624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_69
timestamp 1669390400
transform 1 0 9072 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_550
timestamp 1669390400
transform 1 0 62944 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_554
timestamp 1669390400
transform 1 0 63392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_562
timestamp 1669390400
transform 1 0 64288 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_566
timestamp 1669390400
transform 1 0 64736 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1669390400
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1669390400
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1669390400
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1669390400
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1669390400
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1669390400
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1669390400
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1669390400
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1669390400
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1669390400
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1669390400
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1669390400
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1669390400
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1669390400
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_996
timestamp 1669390400
transform 1 0 112896 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1004
timestamp 1669390400
transform 1 0 113792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1008
timestamp 1669390400
transform 1 0 114240 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_1011
timestamp 1669390400
transform 1 0 114576 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_1027
timestamp 1669390400
transform 1 0 116368 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1029
timestamp 1669390400
transform 1 0 116592 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_1032
timestamp 1669390400
transform 1 0 116928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1040
timestamp 1669390400
transform 1 0 117824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1044
timestamp 1669390400
transform 1 0 118272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_19
timestamp 1669390400
transform 1 0 3472 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_409
timestamp 1669390400
transform 1 0 47152 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_413
timestamp 1669390400
transform 1 0 47600 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_417
timestamp 1669390400
transform 1 0 48048 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_449
timestamp 1669390400
transform 1 0 51632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_457
timestamp 1669390400
transform 1 0 52528 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1669390400
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1669390400
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1669390400
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1669390400
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1669390400
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1669390400
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1669390400
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1669390400
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1669390400
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1669390400
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1669390400
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_960
timestamp 1669390400
transform 1 0 108864 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_992
timestamp 1669390400
transform 1 0 112448 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1008
timestamp 1669390400
transform 1 0 114240 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1012
timestamp 1669390400
transform 1 0 114688 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1027
timestamp 1669390400
transform 1 0 116368 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1031
timestamp 1669390400
transform 1 0 116816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1038
timestamp 1669390400
transform 1 0 117600 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1042
timestamp 1669390400
transform 1 0 118048 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1044
timestamp 1669390400
transform 1 0 118272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_373
timestamp 1669390400
transform 1 0 43120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_381
timestamp 1669390400
transform 1 0 44016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_385
timestamp 1669390400
transform 1 0 44464 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_416
timestamp 1669390400
transform 1 0 47936 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_420
timestamp 1669390400
transform 1 0 48384 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_424
timestamp 1669390400
transform 1 0 48832 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1669390400
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1669390400
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1669390400
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1669390400
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1669390400
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1669390400
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1669390400
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1669390400
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1669390400
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1669390400
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1669390400
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1669390400
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1669390400
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1669390400
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_996
timestamp 1669390400
transform 1 0 112896 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_1028
timestamp 1669390400
transform 1 0 116480 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1044
timestamp 1669390400
transform 1 0 118272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_399
timestamp 1669390400
transform 1 0 46032 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_431
timestamp 1669390400
transform 1 0 49616 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_447
timestamp 1669390400
transform 1 0 51408 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_455
timestamp 1669390400
transform 1 0 52304 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_459
timestamp 1669390400
transform 1 0 52752 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1669390400
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1669390400
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1669390400
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1669390400
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1669390400
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1669390400
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1669390400
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1669390400
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1669390400
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1669390400
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1669390400
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1669390400
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1669390400
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1669390400
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_1031
timestamp 1669390400
transform 1 0 116816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1039
timestamp 1669390400
transform 1 0 117712 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1043
timestamp 1669390400
transform 1 0 118160 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_5
timestamp 1669390400
transform 1 0 1904 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1669390400
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_389
timestamp 1669390400
transform 1 0 44912 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_405
timestamp 1669390400
transform 1 0 46704 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_409
timestamp 1669390400
transform 1 0 47152 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_431
timestamp 1669390400
transform 1 0 49616 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_495
timestamp 1669390400
transform 1 0 56784 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1669390400
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1669390400
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1669390400
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1669390400
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1669390400
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1669390400
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1669390400
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1669390400
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1669390400
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1669390400
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1669390400
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1669390400
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1669390400
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1669390400
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_996
timestamp 1669390400
transform 1 0 112896 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_1028
timestamp 1669390400
transform 1 0 116480 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1044
timestamp 1669390400
transform 1 0 118272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_19
timestamp 1669390400
transform 1 0 3472 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_656
timestamp 1669390400
transform 1 0 74816 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_660
timestamp 1669390400
transform 1 0 75264 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_668
timestamp 1669390400
transform 1 0 76160 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_672
timestamp 1669390400
transform 1 0 76608 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1669390400
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1669390400
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1669390400
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1669390400
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1669390400
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1669390400
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1669390400
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1669390400
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1669390400
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1669390400
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1669390400
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_960
timestamp 1669390400
transform 1 0 108864 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_992
timestamp 1669390400
transform 1 0 112448 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1008
timestamp 1669390400
transform 1 0 114240 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1011
timestamp 1669390400
transform 1 0 114576 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1021
timestamp 1669390400
transform 1 0 115696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1025
timestamp 1669390400
transform 1 0 116144 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1669390400
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1031
timestamp 1669390400
transform 1 0 116816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1038
timestamp 1669390400
transform 1 0 117600 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1042
timestamp 1669390400
transform 1 0 118048 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1044
timestamp 1669390400
transform 1 0 118272 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1669390400
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1669390400
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1669390400
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1669390400
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1669390400
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1669390400
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1669390400
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1669390400
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1669390400
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1669390400
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1669390400
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1669390400
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1669390400
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1669390400
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_996
timestamp 1669390400
transform 1 0 112896 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1012
timestamp 1669390400
transform 1 0 114688 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_1027
timestamp 1669390400
transform 1 0 116368 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_1043
timestamp 1669390400
transform 1 0 118160 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_5
timestamp 1669390400
transform 1 0 1904 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_21
timestamp 1669390400
transform 1 0 3696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_29
timestamp 1669390400
transform 1 0 4592 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_33
timestamp 1669390400
transform 1 0 5040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1669390400
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1669390400
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1669390400
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1669390400
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1669390400
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1669390400
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1669390400
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1669390400
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1669390400
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1669390400
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1669390400
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1669390400
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1669390400
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1669390400
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1669390400
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_1031
timestamp 1669390400
transform 1 0 116816 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1039
timestamp 1669390400
transform 1 0 117712 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_1043
timestamp 1669390400
transform 1 0 118160 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_19
timestamp 1669390400
transform 1 0 3472 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_51
timestamp 1669390400
transform 1 0 7056 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_67
timestamp 1669390400
transform 1 0 8848 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1669390400
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1669390400
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1669390400
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1669390400
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1669390400
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1669390400
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1669390400
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1669390400
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1669390400
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1669390400
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1669390400
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1669390400
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1669390400
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1669390400
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1669390400
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1669390400
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_996
timestamp 1669390400
transform 1 0 112896 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1012
timestamp 1669390400
transform 1 0 114688 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1016
timestamp 1669390400
transform 1 0 115136 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1020
timestamp 1669390400
transform 1 0 115584 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_1037
timestamp 1669390400
transform 1 0 117488 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_5
timestamp 1669390400
transform 1 0 1904 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_21
timestamp 1669390400
transform 1 0 3696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_29
timestamp 1669390400
transform 1 0 4592 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_33
timestamp 1669390400
transform 1 0 5040 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_395
timestamp 1669390400
transform 1 0 45584 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_412
timestamp 1669390400
transform 1 0 47488 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_416
timestamp 1669390400
transform 1 0 47936 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_420
timestamp 1669390400
transform 1 0 48384 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_452
timestamp 1669390400
transform 1 0 51968 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1669390400
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1669390400
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1669390400
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1669390400
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_747
timestamp 1669390400
transform 1 0 85008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_811
timestamp 1669390400
transform 1 0 92176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1669390400
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_818
timestamp 1669390400
transform 1 0 92960 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_882
timestamp 1669390400
transform 1 0 100128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_886
timestamp 1669390400
transform 1 0 100576 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_889
timestamp 1669390400
transform 1 0 100912 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_953
timestamp 1669390400
transform 1 0 108080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_957
timestamp 1669390400
transform 1 0 108528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_960
timestamp 1669390400
transform 1 0 108864 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_992
timestamp 1669390400
transform 1 0 112448 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1008
timestamp 1669390400
transform 1 0 114240 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1012
timestamp 1669390400
transform 1 0 114688 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1027
timestamp 1669390400
transform 1 0 116368 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1031
timestamp 1669390400
transform 1 0 116816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1039
timestamp 1669390400
transform 1 0 117712 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1043
timestamp 1669390400
transform 1 0 118160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_17
timestamp 1669390400
transform 1 0 3248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_21
timestamp 1669390400
transform 1 0 3696 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_53
timestamp 1669390400
transform 1 0 7280 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_69
timestamp 1669390400
transform 1 0 9072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_418
timestamp 1669390400
transform 1 0 48160 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_422
timestamp 1669390400
transform 1 0 48608 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1669390400
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1669390400
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_705
timestamp 1669390400
transform 1 0 80304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1669390400
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_712
timestamp 1669390400
transform 1 0 81088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_776
timestamp 1669390400
transform 1 0 88256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1669390400
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_783
timestamp 1669390400
transform 1 0 89040 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_847
timestamp 1669390400
transform 1 0 96208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1669390400
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_854
timestamp 1669390400
transform 1 0 96992 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_918
timestamp 1669390400
transform 1 0 104160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1669390400
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_925
timestamp 1669390400
transform 1 0 104944 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_989
timestamp 1669390400
transform 1 0 112112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1669390400
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_996
timestamp 1669390400
transform 1 0 112896 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1004
timestamp 1669390400
transform 1 0 113792 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1008
timestamp 1669390400
transform 1 0 114240 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1010
timestamp 1669390400
transform 1 0 114464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1013
timestamp 1669390400
transform 1 0 114800 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1044
timestamp 1669390400
transform 1 0 118272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_19
timestamp 1669390400
transform 1 0 3472 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_394
timestamp 1669390400
transform 1 0 45472 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_401
timestamp 1669390400
transform 1 0 46256 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_433
timestamp 1669390400
transform 1 0 49840 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_449
timestamp 1669390400
transform 1 0 51632 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_457
timestamp 1669390400
transform 1 0 52528 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_495
timestamp 1669390400
transform 1 0 56784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_505
timestamp 1669390400
transform 1 0 57904 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_513
timestamp 1669390400
transform 1 0 58800 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_529
timestamp 1669390400
transform 1 0 60592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1669390400
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1669390400
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1669390400
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_740
timestamp 1669390400
transform 1 0 84224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1669390400
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_747
timestamp 1669390400
transform 1 0 85008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_811
timestamp 1669390400
transform 1 0 92176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1669390400
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_818
timestamp 1669390400
transform 1 0 92960 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_882
timestamp 1669390400
transform 1 0 100128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1669390400
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_889
timestamp 1669390400
transform 1 0 100912 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_953
timestamp 1669390400
transform 1 0 108080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_957
timestamp 1669390400
transform 1 0 108528 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_960
timestamp 1669390400
transform 1 0 108864 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_992
timestamp 1669390400
transform 1 0 112448 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1008
timestamp 1669390400
transform 1 0 114240 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1016
timestamp 1669390400
transform 1 0 115136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1020
timestamp 1669390400
transform 1 0 115584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1669390400
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1031
timestamp 1669390400
transform 1 0 116816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1039
timestamp 1669390400
transform 1 0 117712 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1043
timestamp 1669390400
transform 1 0 118160 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_5
timestamp 1669390400
transform 1 0 1904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_9
timestamp 1669390400
transform 1 0 2352 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_41
timestamp 1669390400
transform 1 0 5936 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_57
timestamp 1669390400
transform 1 0 7728 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_65
timestamp 1669390400
transform 1 0 8624 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_69
timestamp 1669390400
transform 1 0 9072 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1669390400
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1669390400
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_705
timestamp 1669390400
transform 1 0 80304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1669390400
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_712
timestamp 1669390400
transform 1 0 81088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_776
timestamp 1669390400
transform 1 0 88256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1669390400
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_783
timestamp 1669390400
transform 1 0 89040 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_847
timestamp 1669390400
transform 1 0 96208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1669390400
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_854
timestamp 1669390400
transform 1 0 96992 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_918
timestamp 1669390400
transform 1 0 104160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1669390400
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_925
timestamp 1669390400
transform 1 0 104944 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_989
timestamp 1669390400
transform 1 0 112112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_993
timestamp 1669390400
transform 1 0 112560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_996
timestamp 1669390400
transform 1 0 112896 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1004
timestamp 1669390400
transform 1 0 113792 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1008
timestamp 1669390400
transform 1 0 114240 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1011
timestamp 1669390400
transform 1 0 114576 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_1027
timestamp 1669390400
transform 1 0 116368 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1043
timestamp 1669390400
transform 1 0 118160 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_19
timestamp 1669390400
transform 1 0 3472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1669390400
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1669390400
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1669390400
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1669390400
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_669
timestamp 1669390400
transform 1 0 76272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1669390400
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_676
timestamp 1669390400
transform 1 0 77056 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_740
timestamp 1669390400
transform 1 0 84224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_744
timestamp 1669390400
transform 1 0 84672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_747
timestamp 1669390400
transform 1 0 85008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_811
timestamp 1669390400
transform 1 0 92176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_815
timestamp 1669390400
transform 1 0 92624 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_818
timestamp 1669390400
transform 1 0 92960 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_882
timestamp 1669390400
transform 1 0 100128 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_886
timestamp 1669390400
transform 1 0 100576 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_889
timestamp 1669390400
transform 1 0 100912 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_953
timestamp 1669390400
transform 1 0 108080 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_957
timestamp 1669390400
transform 1 0 108528 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_960
timestamp 1669390400
transform 1 0 108864 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_992
timestamp 1669390400
transform 1 0 112448 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1008
timestamp 1669390400
transform 1 0 114240 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1028
timestamp 1669390400
transform 1 0 116480 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1031
timestamp 1669390400
transform 1 0 116816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_1034
timestamp 1669390400
transform 1 0 117152 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1042
timestamp 1669390400
transform 1 0 118048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1044
timestamp 1669390400
transform 1 0 118272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_19
timestamp 1669390400
transform 1 0 3472 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_51
timestamp 1669390400
transform 1 0 7056 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_67
timestamp 1669390400
transform 1 0 8848 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_460
timestamp 1669390400
transform 1 0 52864 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_464
timestamp 1669390400
transform 1 0 53312 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_468
timestamp 1669390400
transform 1 0 53760 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_485
timestamp 1669390400
transform 1 0 55664 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_489
timestamp 1669390400
transform 1 0 56112 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_493
timestamp 1669390400
transform 1 0 56560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_531
timestamp 1669390400
transform 1 0 60816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_535
timestamp 1669390400
transform 1 0 61264 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_542
timestamp 1669390400
transform 1 0 62048 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_558
timestamp 1669390400
transform 1 0 63840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_566
timestamp 1669390400
transform 1 0 64736 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1669390400
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1669390400
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1669390400
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_641
timestamp 1669390400
transform 1 0 73136 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_705
timestamp 1669390400
transform 1 0 80304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_709
timestamp 1669390400
transform 1 0 80752 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_712
timestamp 1669390400
transform 1 0 81088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_776
timestamp 1669390400
transform 1 0 88256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_780
timestamp 1669390400
transform 1 0 88704 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_783
timestamp 1669390400
transform 1 0 89040 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_847
timestamp 1669390400
transform 1 0 96208 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_851
timestamp 1669390400
transform 1 0 96656 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_854
timestamp 1669390400
transform 1 0 96992 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_918
timestamp 1669390400
transform 1 0 104160 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_922
timestamp 1669390400
transform 1 0 104608 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_925
timestamp 1669390400
transform 1 0 104944 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_989
timestamp 1669390400
transform 1 0 112112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_993
timestamp 1669390400
transform 1 0 112560 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_996
timestamp 1669390400
transform 1 0 112896 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_1028
timestamp 1669390400
transform 1 0 116480 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1044
timestamp 1669390400
transform 1 0 118272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_17
timestamp 1669390400
transform 1 0 3248 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_21
timestamp 1669390400
transform 1 0 3696 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_29
timestamp 1669390400
transform 1 0 4592 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_33
timestamp 1669390400
transform 1 0 5040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_493
timestamp 1669390400
transform 1 0 56560 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_525
timestamp 1669390400
transform 1 0 60144 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1669390400
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_564
timestamp 1669390400
transform 1 0 64512 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_596
timestamp 1669390400
transform 1 0 68096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_600
timestamp 1669390400
transform 1 0 68544 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1669390400
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1669390400
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_669
timestamp 1669390400
transform 1 0 76272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1669390400
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_676
timestamp 1669390400
transform 1 0 77056 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_740
timestamp 1669390400
transform 1 0 84224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_744
timestamp 1669390400
transform 1 0 84672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_747
timestamp 1669390400
transform 1 0 85008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_811
timestamp 1669390400
transform 1 0 92176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_815
timestamp 1669390400
transform 1 0 92624 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_818
timestamp 1669390400
transform 1 0 92960 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_882
timestamp 1669390400
transform 1 0 100128 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_886
timestamp 1669390400
transform 1 0 100576 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_889
timestamp 1669390400
transform 1 0 100912 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_953
timestamp 1669390400
transform 1 0 108080 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_957
timestamp 1669390400
transform 1 0 108528 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_960
timestamp 1669390400
transform 1 0 108864 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1024
timestamp 1669390400
transform 1 0 116032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1028
timestamp 1669390400
transform 1 0 116480 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_1031
timestamp 1669390400
transform 1 0 116816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1039
timestamp 1669390400
transform 1 0 117712 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_1043
timestamp 1669390400
transform 1 0 118160 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_460
timestamp 1669390400
transform 1 0 52864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_470
timestamp 1669390400
transform 1 0 53984 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_486
timestamp 1669390400
transform 1 0 55776 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_494
timestamp 1669390400
transform 1 0 56672 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_531
timestamp 1669390400
transform 1 0 60816 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_535
timestamp 1669390400
transform 1 0 61264 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_552
timestamp 1669390400
transform 1 0 63168 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_556
timestamp 1669390400
transform 1 0 63616 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_560
timestamp 1669390400
transform 1 0 64064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1669390400
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1669390400
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1669390400
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_641
timestamp 1669390400
transform 1 0 73136 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_705
timestamp 1669390400
transform 1 0 80304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_709
timestamp 1669390400
transform 1 0 80752 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_712
timestamp 1669390400
transform 1 0 81088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_776
timestamp 1669390400
transform 1 0 88256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_780
timestamp 1669390400
transform 1 0 88704 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_783
timestamp 1669390400
transform 1 0 89040 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_847
timestamp 1669390400
transform 1 0 96208 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_851
timestamp 1669390400
transform 1 0 96656 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_854
timestamp 1669390400
transform 1 0 96992 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_918
timestamp 1669390400
transform 1 0 104160 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_922
timestamp 1669390400
transform 1 0 104608 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_925
timestamp 1669390400
transform 1 0 104944 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_989
timestamp 1669390400
transform 1 0 112112 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_993
timestamp 1669390400
transform 1 0 112560 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_996
timestamp 1669390400
transform 1 0 112896 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_1028
timestamp 1669390400
transform 1 0 116480 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1036
timestamp 1669390400
transform 1 0 117376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1044
timestamp 1669390400
transform 1 0 118272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_17
timestamp 1669390400
transform 1 0 3248 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_21
timestamp 1669390400
transform 1 0 3696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_29
timestamp 1669390400
transform 1 0 4592 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_33
timestamp 1669390400
transform 1 0 5040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_408
timestamp 1669390400
transform 1 0 47040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_410
timestamp 1669390400
transform 1 0 47264 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_413
timestamp 1669390400
transform 1 0 47600 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_430
timestamp 1669390400
transform 1 0 49504 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_434
timestamp 1669390400
transform 1 0 49952 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_438
timestamp 1669390400
transform 1 0 50400 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_442
timestamp 1669390400
transform 1 0 50848 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_444
timestamp 1669390400
transform 1 0 51072 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_447
timestamp 1669390400
transform 1 0 51408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_455
timestamp 1669390400
transform 1 0 52304 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_459
timestamp 1669390400
transform 1 0 52752 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_466
timestamp 1669390400
transform 1 0 53536 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_530
timestamp 1669390400
transform 1 0 60704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1669390400
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1669390400
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_605
timestamp 1669390400
transform 1 0 69104 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_669
timestamp 1669390400
transform 1 0 76272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1669390400
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_676
timestamp 1669390400
transform 1 0 77056 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_740
timestamp 1669390400
transform 1 0 84224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_744
timestamp 1669390400
transform 1 0 84672 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_747
timestamp 1669390400
transform 1 0 85008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_811
timestamp 1669390400
transform 1 0 92176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_815
timestamp 1669390400
transform 1 0 92624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_818
timestamp 1669390400
transform 1 0 92960 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_882
timestamp 1669390400
transform 1 0 100128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_886
timestamp 1669390400
transform 1 0 100576 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_889
timestamp 1669390400
transform 1 0 100912 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_953
timestamp 1669390400
transform 1 0 108080 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_957
timestamp 1669390400
transform 1 0 108528 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_960
timestamp 1669390400
transform 1 0 108864 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1024
timestamp 1669390400
transform 1 0 116032 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1028
timestamp 1669390400
transform 1 0 116480 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1031
timestamp 1669390400
transform 1 0 116816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_1034
timestamp 1669390400
transform 1 0 117152 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_1042
timestamp 1669390400
transform 1 0 118048 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1044
timestamp 1669390400
transform 1 0 118272 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_5
timestamp 1669390400
transform 1 0 1904 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_69
timestamp 1669390400
transform 1 0 9072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_389
timestamp 1669390400
transform 1 0 44912 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_393
timestamp 1669390400
transform 1 0 45360 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_395
timestamp 1669390400
transform 1 0 45584 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_431
timestamp 1669390400
transform 1 0 49616 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_445
timestamp 1669390400
transform 1 0 51184 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_449
timestamp 1669390400
transform 1 0 51632 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_453
timestamp 1669390400
transform 1 0 52080 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_456
timestamp 1669390400
transform 1 0 52416 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_460
timestamp 1669390400
transform 1 0 52864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_464
timestamp 1669390400
transform 1 0 53312 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_468
timestamp 1669390400
transform 1 0 53760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_472
timestamp 1669390400
transform 1 0 54208 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_476
timestamp 1669390400
transform 1 0 54656 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_531
timestamp 1669390400
transform 1 0 60816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_539
timestamp 1669390400
transform 1 0 61712 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_543
timestamp 1669390400
transform 1 0 62160 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_547
timestamp 1669390400
transform 1 0 62608 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1669390400
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1669390400
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1669390400
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1669390400
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1669390400
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_641
timestamp 1669390400
transform 1 0 73136 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_705
timestamp 1669390400
transform 1 0 80304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_709
timestamp 1669390400
transform 1 0 80752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_712
timestamp 1669390400
transform 1 0 81088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_776
timestamp 1669390400
transform 1 0 88256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_780
timestamp 1669390400
transform 1 0 88704 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_783
timestamp 1669390400
transform 1 0 89040 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_847
timestamp 1669390400
transform 1 0 96208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_851
timestamp 1669390400
transform 1 0 96656 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_854
timestamp 1669390400
transform 1 0 96992 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_918
timestamp 1669390400
transform 1 0 104160 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_922
timestamp 1669390400
transform 1 0 104608 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_925
timestamp 1669390400
transform 1 0 104944 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_989
timestamp 1669390400
transform 1 0 112112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_993
timestamp 1669390400
transform 1 0 112560 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_996
timestamp 1669390400
transform 1 0 112896 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1012
timestamp 1669390400
transform 1 0 114688 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_1029
timestamp 1669390400
transform 1 0 116592 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1031
timestamp 1669390400
transform 1 0 116816 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1038
timestamp 1669390400
transform 1 0 117600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_1042
timestamp 1669390400
transform 1 0 118048 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1044
timestamp 1669390400
transform 1 0 118272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_19
timestamp 1669390400
transform 1 0 3472 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_408
timestamp 1669390400
transform 1 0 47040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_416
timestamp 1669390400
transform 1 0 47936 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_424
timestamp 1669390400
transform 1 0 48832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_426
timestamp 1669390400
transform 1 0 49056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_429
timestamp 1669390400
transform 1 0 49392 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_493
timestamp 1669390400
transform 1 0 56560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_497
timestamp 1669390400
transform 1 0 57008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_500
timestamp 1669390400
transform 1 0 57344 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_504
timestamp 1669390400
transform 1 0 57792 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_506
timestamp 1669390400
transform 1 0 58016 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_509
timestamp 1669390400
transform 1 0 58352 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_513
timestamp 1669390400
transform 1 0 58800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_517
timestamp 1669390400
transform 1 0 59248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_521
timestamp 1669390400
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_527
timestamp 1669390400
transform 1 0 60368 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1669390400
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_541
timestamp 1669390400
transform 1 0 61936 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_545
timestamp 1669390400
transform 1 0 62384 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_549
timestamp 1669390400
transform 1 0 62832 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_581
timestamp 1669390400
transform 1 0 66416 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_597
timestamp 1669390400
transform 1 0 68208 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_601
timestamp 1669390400
transform 1 0 68656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1669390400
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_669
timestamp 1669390400
transform 1 0 76272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1669390400
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_676
timestamp 1669390400
transform 1 0 77056 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_740
timestamp 1669390400
transform 1 0 84224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_744
timestamp 1669390400
transform 1 0 84672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_747
timestamp 1669390400
transform 1 0 85008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_811
timestamp 1669390400
transform 1 0 92176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_815
timestamp 1669390400
transform 1 0 92624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_818
timestamp 1669390400
transform 1 0 92960 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_882
timestamp 1669390400
transform 1 0 100128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_886
timestamp 1669390400
transform 1 0 100576 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_889
timestamp 1669390400
transform 1 0 100912 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_953
timestamp 1669390400
transform 1 0 108080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_957
timestamp 1669390400
transform 1 0 108528 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_960
timestamp 1669390400
transform 1 0 108864 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_992
timestamp 1669390400
transform 1 0 112448 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1008
timestamp 1669390400
transform 1 0 114240 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1012
timestamp 1669390400
transform 1 0 114688 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_1027
timestamp 1669390400
transform 1 0 116368 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1031
timestamp 1669390400
transform 1 0 116816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_1034
timestamp 1669390400
transform 1 0 117152 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_1042
timestamp 1669390400
transform 1 0 118048 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1044
timestamp 1669390400
transform 1 0 118272 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1669390400
transform 1 0 44912 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1669390400
transform 1 0 46704 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1669390400
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1669390400
transform 1 0 48048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_421
timestamp 1669390400
transform 1 0 48496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_479
timestamp 1669390400
transform 1 0 54992 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_483
timestamp 1669390400
transform 1 0 55440 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_487
timestamp 1669390400
transform 1 0 55888 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_491
timestamp 1669390400
transform 1 0 56336 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_493
timestamp 1669390400
transform 1 0 56560 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_502
timestamp 1669390400
transform 1 0 57568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_510
timestamp 1669390400
transform 1 0 58464 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_525
timestamp 1669390400
transform 1 0 60144 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_529
timestamp 1669390400
transform 1 0 60592 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_562
timestamp 1669390400
transform 1 0 64288 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_566
timestamp 1669390400
transform 1 0 64736 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1669390400
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1669390400
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1669390400
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_641
timestamp 1669390400
transform 1 0 73136 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_705
timestamp 1669390400
transform 1 0 80304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_709
timestamp 1669390400
transform 1 0 80752 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_712
timestamp 1669390400
transform 1 0 81088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_776
timestamp 1669390400
transform 1 0 88256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_780
timestamp 1669390400
transform 1 0 88704 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_783
timestamp 1669390400
transform 1 0 89040 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_847
timestamp 1669390400
transform 1 0 96208 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_851
timestamp 1669390400
transform 1 0 96656 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_854
timestamp 1669390400
transform 1 0 96992 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_918
timestamp 1669390400
transform 1 0 104160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_922
timestamp 1669390400
transform 1 0 104608 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_925
timestamp 1669390400
transform 1 0 104944 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_989
timestamp 1669390400
transform 1 0 112112 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_993
timestamp 1669390400
transform 1 0 112560 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_996
timestamp 1669390400
transform 1 0 112896 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1004
timestamp 1669390400
transform 1 0 113792 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1008
timestamp 1669390400
transform 1 0 114240 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_1011
timestamp 1669390400
transform 1 0 114576 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_1027
timestamp 1669390400
transform 1 0 116368 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_1043
timestamp 1669390400
transform 1 0 118160 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_408
timestamp 1669390400
transform 1 0 47040 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_412
timestamp 1669390400
transform 1 0 47488 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_415
timestamp 1669390400
transform 1 0 47824 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_419
timestamp 1669390400
transform 1 0 48272 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_427
timestamp 1669390400
transform 1 0 49168 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_443
timestamp 1669390400
transform 1 0 50960 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_459
timestamp 1669390400
transform 1 0 52752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_470
timestamp 1669390400
transform 1 0 53984 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_474
timestamp 1669390400
transform 1 0 54432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_480
timestamp 1669390400
transform 1 0 55104 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_484
timestamp 1669390400
transform 1 0 55552 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_488
timestamp 1669390400
transform 1 0 56000 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_492
timestamp 1669390400
transform 1 0 56448 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_496
timestamp 1669390400
transform 1 0 56896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_500
timestamp 1669390400
transform 1 0 57344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_511
timestamp 1669390400
transform 1 0 58576 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_527
timestamp 1669390400
transform 1 0 60368 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1669390400
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_541
timestamp 1669390400
transform 1 0 61936 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_545
timestamp 1669390400
transform 1 0 62384 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_549
timestamp 1669390400
transform 1 0 62832 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_553
timestamp 1669390400
transform 1 0 63280 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_557
timestamp 1669390400
transform 1 0 63728 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_561
timestamp 1669390400
transform 1 0 64176 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_565
timestamp 1669390400
transform 1 0 64624 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_597
timestamp 1669390400
transform 1 0 68208 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_601
timestamp 1669390400
transform 1 0 68656 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1669390400
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_669
timestamp 1669390400
transform 1 0 76272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1669390400
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_676
timestamp 1669390400
transform 1 0 77056 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_740
timestamp 1669390400
transform 1 0 84224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_744
timestamp 1669390400
transform 1 0 84672 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_747
timestamp 1669390400
transform 1 0 85008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_811
timestamp 1669390400
transform 1 0 92176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_815
timestamp 1669390400
transform 1 0 92624 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_818
timestamp 1669390400
transform 1 0 92960 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_882
timestamp 1669390400
transform 1 0 100128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_886
timestamp 1669390400
transform 1 0 100576 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_889
timestamp 1669390400
transform 1 0 100912 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_953
timestamp 1669390400
transform 1 0 108080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_957
timestamp 1669390400
transform 1 0 108528 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_960
timestamp 1669390400
transform 1 0 108864 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1024
timestamp 1669390400
transform 1 0 116032 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1028
timestamp 1669390400
transform 1 0 116480 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_1031
timestamp 1669390400
transform 1 0 116816 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1039
timestamp 1669390400
transform 1 0 117712 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_1043
timestamp 1669390400
transform 1 0 118160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1669390400
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1669390400
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1669390400
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_421
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_444
timestamp 1669390400
transform 1 0 51072 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_458
timestamp 1669390400
transform 1 0 52640 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_462
timestamp 1669390400
transform 1 0 53088 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_493
timestamp 1669390400
transform 1 0 56560 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_503
timestamp 1669390400
transform 1 0 57680 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_517
timestamp 1669390400
transform 1 0 59248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_531
timestamp 1669390400
transform 1 0 60816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_535
timestamp 1669390400
transform 1 0 61264 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_549
timestamp 1669390400
transform 1 0 62832 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_553
timestamp 1669390400
transform 1 0 63280 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_557
timestamp 1669390400
transform 1 0 63728 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_561
timestamp 1669390400
transform 1 0 64176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_565
timestamp 1669390400
transform 1 0 64624 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1669390400
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_570
timestamp 1669390400
transform 1 0 65184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_573
timestamp 1669390400
transform 1 0 65520 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_577
timestamp 1669390400
transform 1 0 65968 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_580
timestamp 1669390400
transform 1 0 66304 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_598
timestamp 1669390400
transform 1 0 68320 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_630
timestamp 1669390400
transform 1 0 71904 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1669390400
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_641
timestamp 1669390400
transform 1 0 73136 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_705
timestamp 1669390400
transform 1 0 80304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_709
timestamp 1669390400
transform 1 0 80752 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_712
timestamp 1669390400
transform 1 0 81088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_716
timestamp 1669390400
transform 1 0 81536 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_718
timestamp 1669390400
transform 1 0 81760 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_769
timestamp 1669390400
transform 1 0 87472 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_773
timestamp 1669390400
transform 1 0 87920 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_783
timestamp 1669390400
transform 1 0 89040 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_847
timestamp 1669390400
transform 1 0 96208 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_851
timestamp 1669390400
transform 1 0 96656 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_854
timestamp 1669390400
transform 1 0 96992 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_918
timestamp 1669390400
transform 1 0 104160 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_922
timestamp 1669390400
transform 1 0 104608 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_925
timestamp 1669390400
transform 1 0 104944 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_989
timestamp 1669390400
transform 1 0 112112 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_993
timestamp 1669390400
transform 1 0 112560 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_996
timestamp 1669390400
transform 1 0 112896 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1012
timestamp 1669390400
transform 1 0 114688 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_1029
timestamp 1669390400
transform 1 0 116592 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_1033
timestamp 1669390400
transform 1 0 117040 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1041
timestamp 1669390400
transform 1 0 117936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1669390400
transform 1 0 47040 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_416
timestamp 1669390400
transform 1 0 47936 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_419
timestamp 1669390400
transform 1 0 48272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_423
timestamp 1669390400
transform 1 0 48720 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_425
timestamp 1669390400
transform 1 0 48944 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_428
timestamp 1669390400
transform 1 0 49280 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_432
timestamp 1669390400
transform 1 0 49728 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_436
timestamp 1669390400
transform 1 0 50176 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_440
timestamp 1669390400
transform 1 0 50624 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_444
timestamp 1669390400
transform 1 0 51072 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_448
timestamp 1669390400
transform 1 0 51520 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_458
timestamp 1669390400
transform 1 0 52640 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_474
timestamp 1669390400
transform 1 0 54432 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_484
timestamp 1669390400
transform 1 0 55552 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_486
timestamp 1669390400
transform 1 0 55776 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_489
timestamp 1669390400
transform 1 0 56112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_495
timestamp 1669390400
transform 1 0 56784 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_528
timestamp 1669390400
transform 1 0 60480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_542
timestamp 1669390400
transform 1 0 62048 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_576
timestamp 1669390400
transform 1 0 65856 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_580
timestamp 1669390400
transform 1 0 66304 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_582
timestamp 1669390400
transform 1 0 66528 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_592
timestamp 1669390400
transform 1 0 67648 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_596
timestamp 1669390400
transform 1 0 68096 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_600
timestamp 1669390400
transform 1 0 68544 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1669390400
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1669390400
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_669
timestamp 1669390400
transform 1 0 76272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1669390400
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_676
timestamp 1669390400
transform 1 0 77056 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_740
timestamp 1669390400
transform 1 0 84224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_744
timestamp 1669390400
transform 1 0 84672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_747
timestamp 1669390400
transform 1 0 85008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_811
timestamp 1669390400
transform 1 0 92176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_815
timestamp 1669390400
transform 1 0 92624 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_818
timestamp 1669390400
transform 1 0 92960 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_882
timestamp 1669390400
transform 1 0 100128 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_886
timestamp 1669390400
transform 1 0 100576 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_889
timestamp 1669390400
transform 1 0 100912 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_953
timestamp 1669390400
transform 1 0 108080 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_957
timestamp 1669390400
transform 1 0 108528 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_960
timestamp 1669390400
transform 1 0 108864 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1024
timestamp 1669390400
transform 1 0 116032 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1028
timestamp 1669390400
transform 1 0 116480 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_1031
timestamp 1669390400
transform 1 0 116816 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1039
timestamp 1669390400
transform 1 0 117712 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_1043
timestamp 1669390400
transform 1 0 118160 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_361
timestamp 1669390400
transform 1 0 41776 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_369
timestamp 1669390400
transform 1 0 42672 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_373
timestamp 1669390400
transform 1 0 43120 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_405
timestamp 1669390400
transform 1 0 46704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_409
timestamp 1669390400
transform 1 0 47152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_417
timestamp 1669390400
transform 1 0 48048 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_424
timestamp 1669390400
transform 1 0 48832 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_431
timestamp 1669390400
transform 1 0 49616 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_441
timestamp 1669390400
transform 1 0 50736 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_445
timestamp 1669390400
transform 1 0 51184 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_449
timestamp 1669390400
transform 1 0 51632 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_453
timestamp 1669390400
transform 1 0 52080 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_457
timestamp 1669390400
transform 1 0 52528 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_461
timestamp 1669390400
transform 1 0 52976 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_464
timestamp 1669390400
transform 1 0 53312 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_468
timestamp 1669390400
transform 1 0 53760 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_472
timestamp 1669390400
transform 1 0 54208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_476
timestamp 1669390400
transform 1 0 54656 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_480
timestamp 1669390400
transform 1 0 55104 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_484
timestamp 1669390400
transform 1 0 55552 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_488
timestamp 1669390400
transform 1 0 56000 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_502
timestamp 1669390400
transform 1 0 57568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_506
timestamp 1669390400
transform 1 0 58016 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_515
timestamp 1669390400
transform 1 0 59024 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_522
timestamp 1669390400
transform 1 0 59808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_526
timestamp 1669390400
transform 1 0 60256 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_530
timestamp 1669390400
transform 1 0 60704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_534
timestamp 1669390400
transform 1 0 61152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_536
timestamp 1669390400
transform 1 0 61376 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_539
timestamp 1669390400
transform 1 0 61712 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_543
timestamp 1669390400
transform 1 0 62160 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_558
timestamp 1669390400
transform 1 0 63840 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_562
timestamp 1669390400
transform 1 0 64288 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_566
timestamp 1669390400
transform 1 0 64736 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_570
timestamp 1669390400
transform 1 0 65184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_573
timestamp 1669390400
transform 1 0 65520 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_577
timestamp 1669390400
transform 1 0 65968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_583
timestamp 1669390400
transform 1 0 66640 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_587
timestamp 1669390400
transform 1 0 67088 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_619
timestamp 1669390400
transform 1 0 70672 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_635
timestamp 1669390400
transform 1 0 72464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_641
timestamp 1669390400
transform 1 0 73136 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_705
timestamp 1669390400
transform 1 0 80304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_709
timestamp 1669390400
transform 1 0 80752 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_712
timestamp 1669390400
transform 1 0 81088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_776
timestamp 1669390400
transform 1 0 88256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_780
timestamp 1669390400
transform 1 0 88704 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_783
timestamp 1669390400
transform 1 0 89040 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_847
timestamp 1669390400
transform 1 0 96208 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_851
timestamp 1669390400
transform 1 0 96656 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_854
timestamp 1669390400
transform 1 0 96992 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_918
timestamp 1669390400
transform 1 0 104160 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_922
timestamp 1669390400
transform 1 0 104608 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_925
timestamp 1669390400
transform 1 0 104944 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_989
timestamp 1669390400
transform 1 0 112112 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_993
timestamp 1669390400
transform 1 0 112560 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_996
timestamp 1669390400
transform 1 0 112896 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_1030
timestamp 1669390400
transform 1 0 116704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1038
timestamp 1669390400
transform 1 0 117600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_1042
timestamp 1669390400
transform 1 0 118048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1044
timestamp 1669390400
transform 1 0 118272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_17
timestamp 1669390400
transform 1 0 3248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_21
timestamp 1669390400
transform 1 0 3696 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1669390400
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1669390400
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_423
timestamp 1669390400
transform 1 0 48720 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_429
timestamp 1669390400
transform 1 0 49392 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_433
timestamp 1669390400
transform 1 0 49840 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_437
timestamp 1669390400
transform 1 0 50288 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_445
timestamp 1669390400
transform 1 0 51184 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_447
timestamp 1669390400
transform 1 0 51408 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_450
timestamp 1669390400
transform 1 0 51744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_465
timestamp 1669390400
transform 1 0 53424 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_468
timestamp 1669390400
transform 1 0 53760 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_472
timestamp 1669390400
transform 1 0 54208 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_505
timestamp 1669390400
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_509
timestamp 1669390400
transform 1 0 58352 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_515
timestamp 1669390400
transform 1 0 59024 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_519
timestamp 1669390400
transform 1 0 59472 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_522
timestamp 1669390400
transform 1 0 59808 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_526
timestamp 1669390400
transform 1 0 60256 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_530
timestamp 1669390400
transform 1 0 60704 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_585
timestamp 1669390400
transform 1 0 66864 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_589
timestamp 1669390400
transform 1 0 67312 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_593
timestamp 1669390400
transform 1 0 67760 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_597
timestamp 1669390400
transform 1 0 68208 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_601
timestamp 1669390400
transform 1 0 68656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_605
timestamp 1669390400
transform 1 0 69104 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_669
timestamp 1669390400
transform 1 0 76272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1669390400
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_676
timestamp 1669390400
transform 1 0 77056 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_740
timestamp 1669390400
transform 1 0 84224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_744
timestamp 1669390400
transform 1 0 84672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_747
timestamp 1669390400
transform 1 0 85008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_811
timestamp 1669390400
transform 1 0 92176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_815
timestamp 1669390400
transform 1 0 92624 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_818
timestamp 1669390400
transform 1 0 92960 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_882
timestamp 1669390400
transform 1 0 100128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_886
timestamp 1669390400
transform 1 0 100576 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_889
timestamp 1669390400
transform 1 0 100912 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_953
timestamp 1669390400
transform 1 0 108080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_957
timestamp 1669390400
transform 1 0 108528 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_960
timestamp 1669390400
transform 1 0 108864 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_992
timestamp 1669390400
transform 1 0 112448 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1008
timestamp 1669390400
transform 1 0 114240 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1012
timestamp 1669390400
transform 1 0 114688 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_1027
timestamp 1669390400
transform 1 0 116368 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_1031
timestamp 1669390400
transform 1 0 116816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1039
timestamp 1669390400
transform 1 0 117712 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_1043
timestamp 1669390400
transform 1 0 118160 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_17
timestamp 1669390400
transform 1 0 3248 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_49
timestamp 1669390400
transform 1 0 6832 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_65
timestamp 1669390400
transform 1 0 8624 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_69
timestamp 1669390400
transform 1 0 9072 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_389
timestamp 1669390400
transform 1 0 44912 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_407
timestamp 1669390400
transform 1 0 46928 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_417
timestamp 1669390400
transform 1 0 48048 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_436
timestamp 1669390400
transform 1 0 50176 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_467
timestamp 1669390400
transform 1 0 53648 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_471
timestamp 1669390400
transform 1 0 54096 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_474
timestamp 1669390400
transform 1 0 54432 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_478
timestamp 1669390400
transform 1 0 54880 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_482
timestamp 1669390400
transform 1 0 55328 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_490
timestamp 1669390400
transform 1 0 56224 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_494
timestamp 1669390400
transform 1 0 56672 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_502
timestamp 1669390400
transform 1 0 57568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_506
timestamp 1669390400
transform 1 0 58016 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_509
timestamp 1669390400
transform 1 0 58352 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_513
timestamp 1669390400
transform 1 0 58800 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_544
timestamp 1669390400
transform 1 0 62272 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_555
timestamp 1669390400
transform 1 0 63504 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_565
timestamp 1669390400
transform 1 0 64624 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1669390400
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_570
timestamp 1669390400
transform 1 0 65184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_573
timestamp 1669390400
transform 1 0 65520 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_577
timestamp 1669390400
transform 1 0 65968 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_581
timestamp 1669390400
transform 1 0 66416 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_585
timestamp 1669390400
transform 1 0 66864 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_589
timestamp 1669390400
transform 1 0 67312 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_624
timestamp 1669390400
transform 1 0 71232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_632
timestamp 1669390400
transform 1 0 72128 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_636
timestamp 1669390400
transform 1 0 72576 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1669390400
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_641
timestamp 1669390400
transform 1 0 73136 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_705
timestamp 1669390400
transform 1 0 80304 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_709
timestamp 1669390400
transform 1 0 80752 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_712
timestamp 1669390400
transform 1 0 81088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_776
timestamp 1669390400
transform 1 0 88256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_780
timestamp 1669390400
transform 1 0 88704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_783
timestamp 1669390400
transform 1 0 89040 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_847
timestamp 1669390400
transform 1 0 96208 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_851
timestamp 1669390400
transform 1 0 96656 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_854
timestamp 1669390400
transform 1 0 96992 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_918
timestamp 1669390400
transform 1 0 104160 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_922
timestamp 1669390400
transform 1 0 104608 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_925
timestamp 1669390400
transform 1 0 104944 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_989
timestamp 1669390400
transform 1 0 112112 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_993
timestamp 1669390400
transform 1 0 112560 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_996
timestamp 1669390400
transform 1 0 112896 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_1028
timestamp 1669390400
transform 1 0 116480 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1036
timestamp 1669390400
transform 1 0 117376 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1044
timestamp 1669390400
transform 1 0 118272 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_6
timestamp 1669390400
transform 1 0 2016 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_8
timestamp 1669390400
transform 1 0 2240 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_15
timestamp 1669390400
transform 1 0 3024 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_19
timestamp 1669390400
transform 1 0 3472 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_422
timestamp 1669390400
transform 1 0 48608 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_453
timestamp 1669390400
transform 1 0 52080 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_457
timestamp 1669390400
transform 1 0 52528 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_465
timestamp 1669390400
transform 1 0 53424 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_472
timestamp 1669390400
transform 1 0 54208 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_474
timestamp 1669390400
transform 1 0 54432 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_477
timestamp 1669390400
transform 1 0 54768 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_481
timestamp 1669390400
transform 1 0 55216 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_494
timestamp 1669390400
transform 1 0 56672 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_498
timestamp 1669390400
transform 1 0 57120 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_501
timestamp 1669390400
transform 1 0 57456 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_505
timestamp 1669390400
transform 1 0 57904 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_517
timestamp 1669390400
transform 1 0 59248 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_525
timestamp 1669390400
transform 1 0 60144 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_529
timestamp 1669390400
transform 1 0 60592 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1669390400
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_540
timestamp 1669390400
transform 1 0 61824 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_546
timestamp 1669390400
transform 1 0 62496 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_548
timestamp 1669390400
transform 1 0 62720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_555
timestamp 1669390400
transform 1 0 63504 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_588
timestamp 1669390400
transform 1 0 67200 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_596
timestamp 1669390400
transform 1 0 68096 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_600
timestamp 1669390400
transform 1 0 68544 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1669390400
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_605
timestamp 1669390400
transform 1 0 69104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_608
timestamp 1669390400
transform 1 0 69440 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_612
timestamp 1669390400
transform 1 0 69888 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_614
timestamp 1669390400
transform 1 0 70112 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_644
timestamp 1669390400
transform 1 0 73472 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_648
timestamp 1669390400
transform 1 0 73920 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_664
timestamp 1669390400
transform 1 0 75712 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_672
timestamp 1669390400
transform 1 0 76608 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_676
timestamp 1669390400
transform 1 0 77056 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_740
timestamp 1669390400
transform 1 0 84224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_744
timestamp 1669390400
transform 1 0 84672 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_747
timestamp 1669390400
transform 1 0 85008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_811
timestamp 1669390400
transform 1 0 92176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_815
timestamp 1669390400
transform 1 0 92624 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_818
timestamp 1669390400
transform 1 0 92960 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_882
timestamp 1669390400
transform 1 0 100128 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_886
timestamp 1669390400
transform 1 0 100576 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_889
timestamp 1669390400
transform 1 0 100912 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_953
timestamp 1669390400
transform 1 0 108080 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_957
timestamp 1669390400
transform 1 0 108528 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_960
timestamp 1669390400
transform 1 0 108864 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_1024
timestamp 1669390400
transform 1 0 116032 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1028
timestamp 1669390400
transform 1 0 116480 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1031
timestamp 1669390400
transform 1 0 116816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1038
timestamp 1669390400
transform 1 0 117600 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_1042
timestamp 1669390400
transform 1 0 118048 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1044
timestamp 1669390400
transform 1 0 118272 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_389
timestamp 1669390400
transform 1 0 44912 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_391
timestamp 1669390400
transform 1 0 45136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_394
timestamp 1669390400
transform 1 0 45472 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_398
timestamp 1669390400
transform 1 0 45920 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_402
timestamp 1669390400
transform 1 0 46368 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_412
timestamp 1669390400
transform 1 0 47488 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_420
timestamp 1669390400
transform 1 0 48384 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_422
timestamp 1669390400
transform 1 0 48608 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_434
timestamp 1669390400
transform 1 0 49952 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_473
timestamp 1669390400
transform 1 0 54320 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_487
timestamp 1669390400
transform 1 0 55888 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_491
timestamp 1669390400
transform 1 0 56336 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_493
timestamp 1669390400
transform 1 0 56560 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_501
timestamp 1669390400
transform 1 0 57456 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_504
timestamp 1669390400
transform 1 0 57792 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_517
timestamp 1669390400
transform 1 0 59248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_532
timestamp 1669390400
transform 1 0 60928 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_541
timestamp 1669390400
transform 1 0 61936 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_543
timestamp 1669390400
transform 1 0 62160 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_557
timestamp 1669390400
transform 1 0 63728 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_564
timestamp 1669390400
transform 1 0 64512 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_570
timestamp 1669390400
transform 1 0 65184 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_580
timestamp 1669390400
transform 1 0 66304 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_596
timestamp 1669390400
transform 1 0 68096 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_604
timestamp 1669390400
transform 1 0 68992 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_608
timestamp 1669390400
transform 1 0 69440 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_612
timestamp 1669390400
transform 1 0 69888 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_616
timestamp 1669390400
transform 1 0 70336 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_620
timestamp 1669390400
transform 1 0 70784 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_636
timestamp 1669390400
transform 1 0 72576 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1669390400
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_641
timestamp 1669390400
transform 1 0 73136 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_705
timestamp 1669390400
transform 1 0 80304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_709
timestamp 1669390400
transform 1 0 80752 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_712
timestamp 1669390400
transform 1 0 81088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_776
timestamp 1669390400
transform 1 0 88256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_780
timestamp 1669390400
transform 1 0 88704 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_783
timestamp 1669390400
transform 1 0 89040 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_847
timestamp 1669390400
transform 1 0 96208 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_851
timestamp 1669390400
transform 1 0 96656 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_854
timestamp 1669390400
transform 1 0 96992 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_918
timestamp 1669390400
transform 1 0 104160 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_922
timestamp 1669390400
transform 1 0 104608 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_925
timestamp 1669390400
transform 1 0 104944 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_989
timestamp 1669390400
transform 1 0 112112 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_993
timestamp 1669390400
transform 1 0 112560 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_996
timestamp 1669390400
transform 1 0 112896 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1012
timestamp 1669390400
transform 1 0 114688 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1027
timestamp 1669390400
transform 1 0 116368 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1031
timestamp 1669390400
transform 1 0 116816 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1038
timestamp 1669390400
transform 1 0 117600 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_1042
timestamp 1669390400
transform 1 0 118048 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1044
timestamp 1669390400
transform 1 0 118272 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_7
timestamp 1669390400
transform 1 0 2128 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_23
timestamp 1669390400
transform 1 0 3920 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_31
timestamp 1669390400
transform 1 0 4816 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_394
timestamp 1669390400
transform 1 0 45472 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_397
timestamp 1669390400
transform 1 0 45808 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_401
timestamp 1669390400
transform 1 0 46256 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_405
timestamp 1669390400
transform 1 0 46704 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_409
timestamp 1669390400
transform 1 0 47152 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_413
timestamp 1669390400
transform 1 0 47600 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_417
timestamp 1669390400
transform 1 0 48048 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_421
timestamp 1669390400
transform 1 0 48496 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_425
timestamp 1669390400
transform 1 0 48944 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_441
timestamp 1669390400
transform 1 0 50736 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_449
timestamp 1669390400
transform 1 0 51632 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_455
timestamp 1669390400
transform 1 0 52304 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_459
timestamp 1669390400
transform 1 0 52752 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_466
timestamp 1669390400
transform 1 0 53536 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_474
timestamp 1669390400
transform 1 0 54432 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_488
timestamp 1669390400
transform 1 0 56000 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_494
timestamp 1669390400
transform 1 0 56672 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_498
timestamp 1669390400
transform 1 0 57120 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_508
timestamp 1669390400
transform 1 0 58240 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_528
timestamp 1669390400
transform 1 0 60480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_543
timestamp 1669390400
transform 1 0 62160 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_545
timestamp 1669390400
transform 1 0 62384 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_555
timestamp 1669390400
transform 1 0 63504 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_588
timestamp 1669390400
transform 1 0 67200 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_592
timestamp 1669390400
transform 1 0 67648 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_596
timestamp 1669390400
transform 1 0 68096 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_600
timestamp 1669390400
transform 1 0 68544 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1669390400
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_605
timestamp 1669390400
transform 1 0 69104 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_607
timestamp 1669390400
transform 1 0 69328 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_610
timestamp 1669390400
transform 1 0 69664 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_620
timestamp 1669390400
transform 1 0 70784 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_624
timestamp 1669390400
transform 1 0 71232 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_630
timestamp 1669390400
transform 1 0 71904 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_662
timestamp 1669390400
transform 1 0 75488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_670
timestamp 1669390400
transform 1 0 76384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_676
timestamp 1669390400
transform 1 0 77056 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_740
timestamp 1669390400
transform 1 0 84224 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_744
timestamp 1669390400
transform 1 0 84672 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_747
timestamp 1669390400
transform 1 0 85008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_811
timestamp 1669390400
transform 1 0 92176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_815
timestamp 1669390400
transform 1 0 92624 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_818
timestamp 1669390400
transform 1 0 92960 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_882
timestamp 1669390400
transform 1 0 100128 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_886
timestamp 1669390400
transform 1 0 100576 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_889
timestamp 1669390400
transform 1 0 100912 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_953
timestamp 1669390400
transform 1 0 108080 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_957
timestamp 1669390400
transform 1 0 108528 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_960
timestamp 1669390400
transform 1 0 108864 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_992
timestamp 1669390400
transform 1 0 112448 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1008
timestamp 1669390400
transform 1 0 114240 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1012
timestamp 1669390400
transform 1 0 114688 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_1027
timestamp 1669390400
transform 1 0 116368 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1031
timestamp 1669390400
transform 1 0 116816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_1034
timestamp 1669390400
transform 1 0 117152 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_1042
timestamp 1669390400
transform 1 0 118048 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1044
timestamp 1669390400
transform 1 0 118272 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_391
timestamp 1669390400
transform 1 0 45136 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_395
timestamp 1669390400
transform 1 0 45584 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_399
timestamp 1669390400
transform 1 0 46032 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_403
timestamp 1669390400
transform 1 0 46480 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_413
timestamp 1669390400
transform 1 0 47600 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_417
timestamp 1669390400
transform 1 0 48048 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_432
timestamp 1669390400
transform 1 0 49728 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_444
timestamp 1669390400
transform 1 0 51072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_446
timestamp 1669390400
transform 1 0 51296 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_449
timestamp 1669390400
transform 1 0 51632 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_457
timestamp 1669390400
transform 1 0 52528 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_461
timestamp 1669390400
transform 1 0 52976 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_465
timestamp 1669390400
transform 1 0 53424 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_469
timestamp 1669390400
transform 1 0 53872 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_476
timestamp 1669390400
transform 1 0 54656 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_550
timestamp 1669390400
transform 1 0 62944 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_554
timestamp 1669390400
transform 1 0 63392 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_566
timestamp 1669390400
transform 1 0 64736 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_570
timestamp 1669390400
transform 1 0 65184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_573
timestamp 1669390400
transform 1 0 65520 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_577
timestamp 1669390400
transform 1 0 65968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_594
timestamp 1669390400
transform 1 0 67872 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_598
timestamp 1669390400
transform 1 0 68320 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_602
timestamp 1669390400
transform 1 0 68768 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_606
timestamp 1669390400
transform 1 0 69216 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_618
timestamp 1669390400
transform 1 0 70560 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_628
timestamp 1669390400
transform 1 0 71680 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_636
timestamp 1669390400
transform 1 0 72576 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1669390400
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_641
timestamp 1669390400
transform 1 0 73136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_644
timestamp 1669390400
transform 1 0 73472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_708
timestamp 1669390400
transform 1 0 80640 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_712
timestamp 1669390400
transform 1 0 81088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_776
timestamp 1669390400
transform 1 0 88256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_780
timestamp 1669390400
transform 1 0 88704 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_783
timestamp 1669390400
transform 1 0 89040 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_847
timestamp 1669390400
transform 1 0 96208 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_851
timestamp 1669390400
transform 1 0 96656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_854
timestamp 1669390400
transform 1 0 96992 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_918
timestamp 1669390400
transform 1 0 104160 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_922
timestamp 1669390400
transform 1 0 104608 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_925
timestamp 1669390400
transform 1 0 104944 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_989
timestamp 1669390400
transform 1 0 112112 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_993
timestamp 1669390400
transform 1 0 112560 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_996
timestamp 1669390400
transform 1 0 112896 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_1028
timestamp 1669390400
transform 1 0 116480 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_1032
timestamp 1669390400
transform 1 0 116928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1040
timestamp 1669390400
transform 1 0 117824 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1044
timestamp 1669390400
transform 1 0 118272 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_422
timestamp 1669390400
transform 1 0 48608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_426
timestamp 1669390400
transform 1 0 49056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_429
timestamp 1669390400
transform 1 0 49392 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_433
timestamp 1669390400
transform 1 0 49840 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_446
timestamp 1669390400
transform 1 0 51296 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_455
timestamp 1669390400
transform 1 0 52304 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_457
timestamp 1669390400
transform 1 0 52528 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_465
timestamp 1669390400
transform 1 0 53424 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_468
timestamp 1669390400
transform 1 0 53760 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_475
timestamp 1669390400
transform 1 0 54544 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_486
timestamp 1669390400
transform 1 0 55776 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_515
timestamp 1669390400
transform 1 0 59024 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_525
timestamp 1669390400
transform 1 0 60144 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_529
timestamp 1669390400
transform 1 0 60592 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1669390400
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_551
timestamp 1669390400
transform 1 0 63056 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_559
timestamp 1669390400
transform 1 0 63952 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_568
timestamp 1669390400
transform 1 0 64960 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_572
timestamp 1669390400
transform 1 0 65408 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_576
timestamp 1669390400
transform 1 0 65856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_580
timestamp 1669390400
transform 1 0 66304 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_586
timestamp 1669390400
transform 1 0 66976 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_590
timestamp 1669390400
transform 1 0 67424 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_594
timestamp 1669390400
transform 1 0 67872 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_598
timestamp 1669390400
transform 1 0 68320 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1669390400
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_605
timestamp 1669390400
transform 1 0 69104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_635
timestamp 1669390400
transform 1 0 72464 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_639
timestamp 1669390400
transform 1 0 72912 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_671
timestamp 1669390400
transform 1 0 76496 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_673
timestamp 1669390400
transform 1 0 76720 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_676
timestamp 1669390400
transform 1 0 77056 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_740
timestamp 1669390400
transform 1 0 84224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_744
timestamp 1669390400
transform 1 0 84672 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_747
timestamp 1669390400
transform 1 0 85008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_811
timestamp 1669390400
transform 1 0 92176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_815
timestamp 1669390400
transform 1 0 92624 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_818
timestamp 1669390400
transform 1 0 92960 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_882
timestamp 1669390400
transform 1 0 100128 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_886
timestamp 1669390400
transform 1 0 100576 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_889
timestamp 1669390400
transform 1 0 100912 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_953
timestamp 1669390400
transform 1 0 108080 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_957
timestamp 1669390400
transform 1 0 108528 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_960
timestamp 1669390400
transform 1 0 108864 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_992
timestamp 1669390400
transform 1 0 112448 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1008
timestamp 1669390400
transform 1 0 114240 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1012
timestamp 1669390400
transform 1 0 114688 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_1027
timestamp 1669390400
transform 1 0 116368 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1031
timestamp 1669390400
transform 1 0 116816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1038
timestamp 1669390400
transform 1 0 117600 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_1042
timestamp 1669390400
transform 1 0 118048 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1044
timestamp 1669390400
transform 1 0 118272 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_5
timestamp 1669390400
transform 1 0 1904 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_69
timestamp 1669390400
transform 1 0 9072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_389
timestamp 1669390400
transform 1 0 44912 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_392
timestamp 1669390400
transform 1 0 45248 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_396
timestamp 1669390400
transform 1 0 45696 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_400
timestamp 1669390400
transform 1 0 46144 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_404
timestamp 1669390400
transform 1 0 46592 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_408
timestamp 1669390400
transform 1 0 47040 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_416
timestamp 1669390400
transform 1 0 47936 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_422
timestamp 1669390400
transform 1 0 48608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_432
timestamp 1669390400
transform 1 0 49728 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_436
timestamp 1669390400
transform 1 0 50176 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_444
timestamp 1669390400
transform 1 0 51072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_452
timestamp 1669390400
transform 1 0 51968 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_486
timestamp 1669390400
transform 1 0 55776 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_494
timestamp 1669390400
transform 1 0 56672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_509
timestamp 1669390400
transform 1 0 58352 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_516
timestamp 1669390400
transform 1 0 59136 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_520
timestamp 1669390400
transform 1 0 59584 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_524
timestamp 1669390400
transform 1 0 60032 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_556
timestamp 1669390400
transform 1 0 63616 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_566
timestamp 1669390400
transform 1 0 64736 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_570
timestamp 1669390400
transform 1 0 65184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_577
timestamp 1669390400
transform 1 0 65968 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_581
timestamp 1669390400
transform 1 0 66416 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_585
timestamp 1669390400
transform 1 0 66864 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_589
timestamp 1669390400
transform 1 0 67312 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_593
timestamp 1669390400
transform 1 0 67760 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_597
timestamp 1669390400
transform 1 0 68208 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_605
timestamp 1669390400
transform 1 0 69104 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_609
timestamp 1669390400
transform 1 0 69552 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_613
timestamp 1669390400
transform 1 0 70000 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_615
timestamp 1669390400
transform 1 0 70224 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_618
timestamp 1669390400
transform 1 0 70560 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_628
timestamp 1669390400
transform 1 0 71680 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_636
timestamp 1669390400
transform 1 0 72576 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1669390400
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_641
timestamp 1669390400
transform 1 0 73136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_644
timestamp 1669390400
transform 1 0 73472 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_648
timestamp 1669390400
transform 1 0 73920 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_680
timestamp 1669390400
transform 1 0 77504 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_696
timestamp 1669390400
transform 1 0 79296 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_704
timestamp 1669390400
transform 1 0 80192 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_708
timestamp 1669390400
transform 1 0 80640 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_712
timestamp 1669390400
transform 1 0 81088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_776
timestamp 1669390400
transform 1 0 88256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_780
timestamp 1669390400
transform 1 0 88704 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_783
timestamp 1669390400
transform 1 0 89040 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_847
timestamp 1669390400
transform 1 0 96208 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_851
timestamp 1669390400
transform 1 0 96656 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_854
timestamp 1669390400
transform 1 0 96992 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_918
timestamp 1669390400
transform 1 0 104160 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_922
timestamp 1669390400
transform 1 0 104608 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_925
timestamp 1669390400
transform 1 0 104944 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_989
timestamp 1669390400
transform 1 0 112112 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_993
timestamp 1669390400
transform 1 0 112560 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_996
timestamp 1669390400
transform 1 0 112896 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_1028
timestamp 1669390400
transform 1 0 116480 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1044
timestamp 1669390400
transform 1 0 118272 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_19
timestamp 1669390400
transform 1 0 3472 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_396
timestamp 1669390400
transform 1 0 45696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_400
timestamp 1669390400
transform 1 0 46144 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_404
timestamp 1669390400
transform 1 0 46592 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_408
timestamp 1669390400
transform 1 0 47040 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_412
timestamp 1669390400
transform 1 0 47488 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_416
timestamp 1669390400
transform 1 0 47936 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_420
timestamp 1669390400
transform 1 0 48384 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_424
timestamp 1669390400
transform 1 0 48832 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_432
timestamp 1669390400
transform 1 0 49728 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_440
timestamp 1669390400
transform 1 0 50624 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_446
timestamp 1669390400
transform 1 0 51296 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_450
timestamp 1669390400
transform 1 0 51744 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_459
timestamp 1669390400
transform 1 0 52752 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_469
timestamp 1669390400
transform 1 0 53872 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_480
timestamp 1669390400
transform 1 0 55104 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_492
timestamp 1669390400
transform 1 0 56448 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_496
timestamp 1669390400
transform 1 0 56896 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_500
timestamp 1669390400
transform 1 0 57344 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_504
timestamp 1669390400
transform 1 0 57792 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_506
timestamp 1669390400
transform 1 0 58016 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_509
timestamp 1669390400
transform 1 0 58352 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_520
timestamp 1669390400
transform 1 0 59584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_524
timestamp 1669390400
transform 1 0 60032 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1669390400
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_549
timestamp 1669390400
transform 1 0 62832 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_553
timestamp 1669390400
transform 1 0 63280 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_565
timestamp 1669390400
transform 1 0 64624 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_574
timestamp 1669390400
transform 1 0 65632 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_590
timestamp 1669390400
transform 1 0 67424 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_598
timestamp 1669390400
transform 1 0 68320 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_602
timestamp 1669390400
transform 1 0 68768 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_605
timestamp 1669390400
transform 1 0 69104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_608
timestamp 1669390400
transform 1 0 69440 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_612
timestamp 1669390400
transform 1 0 69888 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_616
timestamp 1669390400
transform 1 0 70336 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_646
timestamp 1669390400
transform 1 0 73696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_650
timestamp 1669390400
transform 1 0 74144 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_666
timestamp 1669390400
transform 1 0 75936 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_676
timestamp 1669390400
transform 1 0 77056 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_740
timestamp 1669390400
transform 1 0 84224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_744
timestamp 1669390400
transform 1 0 84672 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_747
timestamp 1669390400
transform 1 0 85008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_811
timestamp 1669390400
transform 1 0 92176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_815
timestamp 1669390400
transform 1 0 92624 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_818
timestamp 1669390400
transform 1 0 92960 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_882
timestamp 1669390400
transform 1 0 100128 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_886
timestamp 1669390400
transform 1 0 100576 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_889
timestamp 1669390400
transform 1 0 100912 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_953
timestamp 1669390400
transform 1 0 108080 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_957
timestamp 1669390400
transform 1 0 108528 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_960
timestamp 1669390400
transform 1 0 108864 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1024
timestamp 1669390400
transform 1 0 116032 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1028
timestamp 1669390400
transform 1 0 116480 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_1031
timestamp 1669390400
transform 1 0 116816 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1039
timestamp 1669390400
transform 1 0 117712 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_1043
timestamp 1669390400
transform 1 0 118160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_293
timestamp 1669390400
transform 1 0 34160 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_297
timestamp 1669390400
transform 1 0 34608 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_329
timestamp 1669390400
transform 1 0 38192 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_345
timestamp 1669390400
transform 1 0 39984 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_353
timestamp 1669390400
transform 1 0 40880 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_361
timestamp 1669390400
transform 1 0 41776 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_365
timestamp 1669390400
transform 1 0 42224 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_369
timestamp 1669390400
transform 1 0 42672 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_377
timestamp 1669390400
transform 1 0 43568 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_393
timestamp 1669390400
transform 1 0 45360 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_442
timestamp 1669390400
transform 1 0 50848 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_448
timestamp 1669390400
transform 1 0 51520 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_452
timestamp 1669390400
transform 1 0 51968 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_456
timestamp 1669390400
transform 1 0 52416 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_460
timestamp 1669390400
transform 1 0 52864 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_464
timestamp 1669390400
transform 1 0 53312 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_472
timestamp 1669390400
transform 1 0 54208 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_480
timestamp 1669390400
transform 1 0 55104 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_514
timestamp 1669390400
transform 1 0 58912 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_522
timestamp 1669390400
transform 1 0 59808 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_526
timestamp 1669390400
transform 1 0 60256 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_530
timestamp 1669390400
transform 1 0 60704 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_534
timestamp 1669390400
transform 1 0 61152 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_538
timestamp 1669390400
transform 1 0 61600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_542
timestamp 1669390400
transform 1 0 62048 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_546
timestamp 1669390400
transform 1 0 62496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_550
timestamp 1669390400
transform 1 0 62944 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_560
timestamp 1669390400
transform 1 0 64064 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_562
timestamp 1669390400
transform 1 0 64288 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_565
timestamp 1669390400
transform 1 0 64624 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1669390400
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_570
timestamp 1669390400
transform 1 0 65184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_573
timestamp 1669390400
transform 1 0 65520 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_583
timestamp 1669390400
transform 1 0 66640 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_587
timestamp 1669390400
transform 1 0 67088 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_591
timestamp 1669390400
transform 1 0 67536 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_623
timestamp 1669390400
transform 1 0 71120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_641
timestamp 1669390400
transform 1 0 73136 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_705
timestamp 1669390400
transform 1 0 80304 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_709
timestamp 1669390400
transform 1 0 80752 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_712
timestamp 1669390400
transform 1 0 81088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_776
timestamp 1669390400
transform 1 0 88256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_780
timestamp 1669390400
transform 1 0 88704 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_783
timestamp 1669390400
transform 1 0 89040 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_847
timestamp 1669390400
transform 1 0 96208 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_851
timestamp 1669390400
transform 1 0 96656 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_854
timestamp 1669390400
transform 1 0 96992 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_918
timestamp 1669390400
transform 1 0 104160 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_922
timestamp 1669390400
transform 1 0 104608 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_925
timestamp 1669390400
transform 1 0 104944 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_989
timestamp 1669390400
transform 1 0 112112 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_993
timestamp 1669390400
transform 1 0 112560 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_996
timestamp 1669390400
transform 1 0 112896 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1012
timestamp 1669390400
transform 1 0 114688 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_1029
timestamp 1669390400
transform 1 0 116592 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_1033
timestamp 1669390400
transform 1 0 117040 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1041
timestamp 1669390400
transform 1 0 117936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_395
timestamp 1669390400
transform 1 0 45584 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_399
timestamp 1669390400
transform 1 0 46032 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_403
timestamp 1669390400
transform 1 0 46480 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_407
timestamp 1669390400
transform 1 0 46928 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_411
timestamp 1669390400
transform 1 0 47376 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_415
timestamp 1669390400
transform 1 0 47824 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_424
timestamp 1669390400
transform 1 0 48832 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_437
timestamp 1669390400
transform 1 0 50288 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_441
timestamp 1669390400
transform 1 0 50736 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_445
timestamp 1669390400
transform 1 0 51184 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_457
timestamp 1669390400
transform 1 0 52528 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_514
timestamp 1669390400
transform 1 0 58912 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_522
timestamp 1669390400
transform 1 0 59808 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_526
timestamp 1669390400
transform 1 0 60256 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_530
timestamp 1669390400
transform 1 0 60704 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_537
timestamp 1669390400
transform 1 0 61488 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_541
timestamp 1669390400
transform 1 0 61936 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_545
timestamp 1669390400
transform 1 0 62384 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_549
timestamp 1669390400
transform 1 0 62832 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_582
timestamp 1669390400
transform 1 0 66528 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_592
timestamp 1669390400
transform 1 0 67648 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_600
timestamp 1669390400
transform 1 0 68544 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1669390400
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_605
timestamp 1669390400
transform 1 0 69104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_608
timestamp 1669390400
transform 1 0 69440 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_618
timestamp 1669390400
transform 1 0 70560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_622
timestamp 1669390400
transform 1 0 71008 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_626
timestamp 1669390400
transform 1 0 71456 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_658
timestamp 1669390400
transform 1 0 75040 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_676
timestamp 1669390400
transform 1 0 77056 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_740
timestamp 1669390400
transform 1 0 84224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_744
timestamp 1669390400
transform 1 0 84672 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_747
timestamp 1669390400
transform 1 0 85008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_811
timestamp 1669390400
transform 1 0 92176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_815
timestamp 1669390400
transform 1 0 92624 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_818
timestamp 1669390400
transform 1 0 92960 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_882
timestamp 1669390400
transform 1 0 100128 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_886
timestamp 1669390400
transform 1 0 100576 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_889
timestamp 1669390400
transform 1 0 100912 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_953
timestamp 1669390400
transform 1 0 108080 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_957
timestamp 1669390400
transform 1 0 108528 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_960
timestamp 1669390400
transform 1 0 108864 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1024
timestamp 1669390400
transform 1 0 116032 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1028
timestamp 1669390400
transform 1 0 116480 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_1031
timestamp 1669390400
transform 1 0 116816 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1039
timestamp 1669390400
transform 1 0 117712 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_1043
timestamp 1669390400
transform 1 0 118160 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_318
timestamp 1669390400
transform 1 0 36960 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_334
timestamp 1669390400
transform 1 0 38752 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_342
timestamp 1669390400
transform 1 0 39648 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_346
timestamp 1669390400
transform 1 0 40096 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_364
timestamp 1669390400
transform 1 0 42112 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_380
timestamp 1669390400
transform 1 0 43904 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_388
timestamp 1669390400
transform 1 0 44800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_392
timestamp 1669390400
transform 1 0 45248 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_394
timestamp 1669390400
transform 1 0 45472 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_397
timestamp 1669390400
transform 1 0 45808 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_401
timestamp 1669390400
transform 1 0 46256 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_405
timestamp 1669390400
transform 1 0 46704 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_409
timestamp 1669390400
transform 1 0 47152 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_413
timestamp 1669390400
transform 1 0 47600 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_417
timestamp 1669390400
transform 1 0 48048 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_437
timestamp 1669390400
transform 1 0 50288 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_443
timestamp 1669390400
transform 1 0 50960 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_447
timestamp 1669390400
transform 1 0 51408 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_457
timestamp 1669390400
transform 1 0 52528 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_463
timestamp 1669390400
transform 1 0 53200 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_467
timestamp 1669390400
transform 1 0 53648 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_470
timestamp 1669390400
transform 1 0 53984 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_484
timestamp 1669390400
transform 1 0 55552 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_488
timestamp 1669390400
transform 1 0 56000 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_512
timestamp 1669390400
transform 1 0 58688 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_520
timestamp 1669390400
transform 1 0 59584 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_553
timestamp 1669390400
transform 1 0 63280 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_561
timestamp 1669390400
transform 1 0 64176 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_565
timestamp 1669390400
transform 1 0 64624 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_567
timestamp 1669390400
transform 1 0 64848 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_570
timestamp 1669390400
transform 1 0 65184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_573
timestamp 1669390400
transform 1 0 65520 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_581
timestamp 1669390400
transform 1 0 66416 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_584
timestamp 1669390400
transform 1 0 66752 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_588
timestamp 1669390400
transform 1 0 67200 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_591
timestamp 1669390400
transform 1 0 67536 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_599
timestamp 1669390400
transform 1 0 68432 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_603
timestamp 1669390400
transform 1 0 68880 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_607
timestamp 1669390400
transform 1 0 69328 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1669390400
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_641
timestamp 1669390400
transform 1 0 73136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_644
timestamp 1669390400
transform 1 0 73472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_708
timestamp 1669390400
transform 1 0 80640 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_712
timestamp 1669390400
transform 1 0 81088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_776
timestamp 1669390400
transform 1 0 88256 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_780
timestamp 1669390400
transform 1 0 88704 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_783
timestamp 1669390400
transform 1 0 89040 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_793
timestamp 1669390400
transform 1 0 90160 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_825
timestamp 1669390400
transform 1 0 93744 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_841
timestamp 1669390400
transform 1 0 95536 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_849
timestamp 1669390400
transform 1 0 96432 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_851
timestamp 1669390400
transform 1 0 96656 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_854
timestamp 1669390400
transform 1 0 96992 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_918
timestamp 1669390400
transform 1 0 104160 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_922
timestamp 1669390400
transform 1 0 104608 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_925
timestamp 1669390400
transform 1 0 104944 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_989
timestamp 1669390400
transform 1 0 112112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_993
timestamp 1669390400
transform 1 0 112560 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_996
timestamp 1669390400
transform 1 0 112896 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_1028
timestamp 1669390400
transform 1 0 116480 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1044
timestamp 1669390400
transform 1 0 118272 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_7
timestamp 1669390400
transform 1 0 2128 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_23
timestamp 1669390400
transform 1 0 3920 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_31
timestamp 1669390400
transform 1 0 4816 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_337
timestamp 1669390400
transform 1 0 39088 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_343
timestamp 1669390400
transform 1 0 39760 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_347
timestamp 1669390400
transform 1 0 40208 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_355
timestamp 1669390400
transform 1 0 41104 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_387
timestamp 1669390400
transform 1 0 44688 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_398
timestamp 1669390400
transform 1 0 45920 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_415
timestamp 1669390400
transform 1 0 47824 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_417
timestamp 1669390400
transform 1 0 48048 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_420
timestamp 1669390400
transform 1 0 48384 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_424
timestamp 1669390400
transform 1 0 48832 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_428
timestamp 1669390400
transform 1 0 49280 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_436
timestamp 1669390400
transform 1 0 50176 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_440
timestamp 1669390400
transform 1 0 50624 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_450
timestamp 1669390400
transform 1 0 51744 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_476
timestamp 1669390400
transform 1 0 54656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_484
timestamp 1669390400
transform 1 0 55552 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_488
timestamp 1669390400
transform 1 0 56000 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_492
timestamp 1669390400
transform 1 0 56448 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_496
timestamp 1669390400
transform 1 0 56896 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_502
timestamp 1669390400
transform 1 0 57568 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_510
timestamp 1669390400
transform 1 0 58464 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_522
timestamp 1669390400
transform 1 0 59808 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_526
timestamp 1669390400
transform 1 0 60256 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_528
timestamp 1669390400
transform 1 0 60480 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1669390400
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_537
timestamp 1669390400
transform 1 0 61488 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_553
timestamp 1669390400
transform 1 0 63280 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_557
timestamp 1669390400
transform 1 0 63728 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_559
timestamp 1669390400
transform 1 0 63952 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_562
timestamp 1669390400
transform 1 0 64288 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_564
timestamp 1669390400
transform 1 0 64512 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_567
timestamp 1669390400
transform 1 0 64848 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_571
timestamp 1669390400
transform 1 0 65296 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_575
timestamp 1669390400
transform 1 0 65744 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_579
timestamp 1669390400
transform 1 0 66192 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_583
timestamp 1669390400
transform 1 0 66640 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_587
timestamp 1669390400
transform 1 0 67088 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_590
timestamp 1669390400
transform 1 0 67424 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_594
timestamp 1669390400
transform 1 0 67872 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_598
timestamp 1669390400
transform 1 0 68320 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1669390400
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_605
timestamp 1669390400
transform 1 0 69104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_620
timestamp 1669390400
transform 1 0 70784 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_624
timestamp 1669390400
transform 1 0 71232 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_628
timestamp 1669390400
transform 1 0 71680 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_632
timestamp 1669390400
transform 1 0 72128 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_664
timestamp 1669390400
transform 1 0 75712 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_672
timestamp 1669390400
transform 1 0 76608 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_676
timestamp 1669390400
transform 1 0 77056 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_740
timestamp 1669390400
transform 1 0 84224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_744
timestamp 1669390400
transform 1 0 84672 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_747
timestamp 1669390400
transform 1 0 85008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_811
timestamp 1669390400
transform 1 0 92176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_815
timestamp 1669390400
transform 1 0 92624 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_818
timestamp 1669390400
transform 1 0 92960 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_882
timestamp 1669390400
transform 1 0 100128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_886
timestamp 1669390400
transform 1 0 100576 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_889
timestamp 1669390400
transform 1 0 100912 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_953
timestamp 1669390400
transform 1 0 108080 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_957
timestamp 1669390400
transform 1 0 108528 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_960
timestamp 1669390400
transform 1 0 108864 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_992
timestamp 1669390400
transform 1 0 112448 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1008
timestamp 1669390400
transform 1 0 114240 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_1011
timestamp 1669390400
transform 1 0 114576 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_1027
timestamp 1669390400
transform 1 0 116368 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_1031
timestamp 1669390400
transform 1 0 116816 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1039
timestamp 1669390400
transform 1 0 117712 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_1043
timestamp 1669390400
transform 1 0 118160 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1669390400
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_373
timestamp 1669390400
transform 1 0 43120 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_381
timestamp 1669390400
transform 1 0 44016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_385
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_417
timestamp 1669390400
transform 1 0 48048 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_421
timestamp 1669390400
transform 1 0 48496 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1669390400
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_441
timestamp 1669390400
transform 1 0 50736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_445
timestamp 1669390400
transform 1 0 51184 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_449
timestamp 1669390400
transform 1 0 51632 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_453
timestamp 1669390400
transform 1 0 52080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_461
timestamp 1669390400
transform 1 0 52976 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_471
timestamp 1669390400
transform 1 0 54096 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_484
timestamp 1669390400
transform 1 0 55552 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_494
timestamp 1669390400
transform 1 0 56672 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_503
timestamp 1669390400
transform 1 0 57680 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_507
timestamp 1669390400
transform 1 0 58128 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_509
timestamp 1669390400
transform 1 0 58352 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_512
timestamp 1669390400
transform 1 0 58688 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_523
timestamp 1669390400
transform 1 0 59920 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_527
timestamp 1669390400
transform 1 0 60368 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_541
timestamp 1669390400
transform 1 0 61936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_547
timestamp 1669390400
transform 1 0 62608 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_551
timestamp 1669390400
transform 1 0 63056 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_553
timestamp 1669390400
transform 1 0 63280 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_560
timestamp 1669390400
transform 1 0 64064 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_564
timestamp 1669390400
transform 1 0 64512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_570
timestamp 1669390400
transform 1 0 65184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_573
timestamp 1669390400
transform 1 0 65520 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_577
timestamp 1669390400
transform 1 0 65968 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_579
timestamp 1669390400
transform 1 0 66192 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_594
timestamp 1669390400
transform 1 0 67872 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_605
timestamp 1669390400
transform 1 0 69104 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_607
timestamp 1669390400
transform 1 0 69328 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_620
timestamp 1669390400
transform 1 0 70784 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_624
timestamp 1669390400
transform 1 0 71232 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_628
timestamp 1669390400
transform 1 0 71680 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_632
timestamp 1669390400
transform 1 0 72128 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_636
timestamp 1669390400
transform 1 0 72576 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1669390400
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_641
timestamp 1669390400
transform 1 0 73136 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_673
timestamp 1669390400
transform 1 0 76720 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_689
timestamp 1669390400
transform 1 0 78512 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_699
timestamp 1669390400
transform 1 0 79632 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_707
timestamp 1669390400
transform 1 0 80528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_709
timestamp 1669390400
transform 1 0 80752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_712
timestamp 1669390400
transform 1 0 81088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_776
timestamp 1669390400
transform 1 0 88256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_780
timestamp 1669390400
transform 1 0 88704 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_783
timestamp 1669390400
transform 1 0 89040 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_847
timestamp 1669390400
transform 1 0 96208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_851
timestamp 1669390400
transform 1 0 96656 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_854
timestamp 1669390400
transform 1 0 96992 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_918
timestamp 1669390400
transform 1 0 104160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_922
timestamp 1669390400
transform 1 0 104608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_925
timestamp 1669390400
transform 1 0 104944 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_989
timestamp 1669390400
transform 1 0 112112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_993
timestamp 1669390400
transform 1 0 112560 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_996
timestamp 1669390400
transform 1 0 112896 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1004
timestamp 1669390400
transform 1 0 113792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1008
timestamp 1669390400
transform 1 0 114240 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_1011
timestamp 1669390400
transform 1 0 114576 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_1027
timestamp 1669390400
transform 1 0 116368 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_1043
timestamp 1669390400
transform 1 0 118160 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_17
timestamp 1669390400
transform 1 0 3248 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_21
timestamp 1669390400
transform 1 0 3696 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_29
timestamp 1669390400
transform 1 0 4592 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_33
timestamp 1669390400
transform 1 0 5040 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1669390400
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1669390400
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1669390400
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1669390400
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1669390400
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1669390400
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_353
timestamp 1669390400
transform 1 0 40880 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_357
timestamp 1669390400
transform 1 0 41328 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_367
timestamp 1669390400
transform 1 0 42448 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_383
timestamp 1669390400
transform 1 0 44240 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_387
timestamp 1669390400
transform 1 0 44688 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_402
timestamp 1669390400
transform 1 0 46368 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_406
timestamp 1669390400
transform 1 0 46816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_409
timestamp 1669390400
transform 1 0 47152 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_413
timestamp 1669390400
transform 1 0 47600 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_417
timestamp 1669390400
transform 1 0 48048 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_450
timestamp 1669390400
transform 1 0 51744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_456
timestamp 1669390400
transform 1 0 52416 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_496
timestamp 1669390400
transform 1 0 56896 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_503
timestamp 1669390400
transform 1 0 57680 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_507
timestamp 1669390400
transform 1 0 58128 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_511
timestamp 1669390400
transform 1 0 58576 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_515
timestamp 1669390400
transform 1 0 59024 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_519
timestamp 1669390400
transform 1 0 59472 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_527
timestamp 1669390400
transform 1 0 60368 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_531
timestamp 1669390400
transform 1 0 60816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_536
timestamp 1669390400
transform 1 0 61376 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_539
timestamp 1669390400
transform 1 0 61712 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_543
timestamp 1669390400
transform 1 0 62160 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_549
timestamp 1669390400
transform 1 0 62832 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_565
timestamp 1669390400
transform 1 0 64624 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_569
timestamp 1669390400
transform 1 0 65072 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_576
timestamp 1669390400
transform 1 0 65856 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_580
timestamp 1669390400
transform 1 0 66304 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_588
timestamp 1669390400
transform 1 0 67200 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_592
timestamp 1669390400
transform 1 0 67648 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_596
timestamp 1669390400
transform 1 0 68096 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1669390400
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_605
timestamp 1669390400
transform 1 0 69104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_608
timestamp 1669390400
transform 1 0 69440 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_612
timestamp 1669390400
transform 1 0 69888 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_642
timestamp 1669390400
transform 1 0 73248 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_646
timestamp 1669390400
transform 1 0 73696 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_662
timestamp 1669390400
transform 1 0 75488 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_670
timestamp 1669390400
transform 1 0 76384 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_676
timestamp 1669390400
transform 1 0 77056 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_740
timestamp 1669390400
transform 1 0 84224 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_744
timestamp 1669390400
transform 1 0 84672 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_747
timestamp 1669390400
transform 1 0 85008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_811
timestamp 1669390400
transform 1 0 92176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_815
timestamp 1669390400
transform 1 0 92624 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_818
timestamp 1669390400
transform 1 0 92960 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_882
timestamp 1669390400
transform 1 0 100128 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_886
timestamp 1669390400
transform 1 0 100576 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_889
timestamp 1669390400
transform 1 0 100912 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_953
timestamp 1669390400
transform 1 0 108080 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_957
timestamp 1669390400
transform 1 0 108528 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_960
timestamp 1669390400
transform 1 0 108864 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1024
timestamp 1669390400
transform 1 0 116032 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1028
timestamp 1669390400
transform 1 0 116480 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_1031
timestamp 1669390400
transform 1 0 116816 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1039
timestamp 1669390400
transform 1 0 117712 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1044
timestamp 1669390400
transform 1 0 118272 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_66
timestamp 1669390400
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1669390400
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1669390400
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1669390400
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1669390400
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1669390400
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1669390400
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1669390400
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_389
timestamp 1669390400
transform 1 0 44912 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_405
timestamp 1669390400
transform 1 0 46704 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_413
timestamp 1669390400
transform 1 0 47600 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_417
timestamp 1669390400
transform 1 0 48048 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_421
timestamp 1669390400
transform 1 0 48496 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1669390400
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_435
timestamp 1669390400
transform 1 0 50064 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_441
timestamp 1669390400
transform 1 0 50736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_445
timestamp 1669390400
transform 1 0 51184 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_449
timestamp 1669390400
transform 1 0 51632 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_453
timestamp 1669390400
transform 1 0 52080 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_457
timestamp 1669390400
transform 1 0 52528 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_467
timestamp 1669390400
transform 1 0 53648 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_471
timestamp 1669390400
transform 1 0 54096 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_474
timestamp 1669390400
transform 1 0 54432 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_478
timestamp 1669390400
transform 1 0 54880 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_482
timestamp 1669390400
transform 1 0 55328 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_486
timestamp 1669390400
transform 1 0 55776 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_490
timestamp 1669390400
transform 1 0 56224 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1669390400
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_537
timestamp 1669390400
transform 1 0 61488 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_547
timestamp 1669390400
transform 1 0 62608 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_551
timestamp 1669390400
transform 1 0 63056 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1669390400
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_570
timestamp 1669390400
transform 1 0 65184 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_572
timestamp 1669390400
transform 1 0 65408 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_602
timestamp 1669390400
transform 1 0 68768 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_612
timestamp 1669390400
transform 1 0 69888 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_621
timestamp 1669390400
transform 1 0 70896 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_625
timestamp 1669390400
transform 1 0 71344 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_629
timestamp 1669390400
transform 1 0 71792 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_637
timestamp 1669390400
transform 1 0 72688 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_641
timestamp 1669390400
transform 1 0 73136 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_705
timestamp 1669390400
transform 1 0 80304 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_709
timestamp 1669390400
transform 1 0 80752 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_712
timestamp 1669390400
transform 1 0 81088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_776
timestamp 1669390400
transform 1 0 88256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_780
timestamp 1669390400
transform 1 0 88704 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_783
timestamp 1669390400
transform 1 0 89040 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_847
timestamp 1669390400
transform 1 0 96208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_851
timestamp 1669390400
transform 1 0 96656 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_854
timestamp 1669390400
transform 1 0 96992 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_918
timestamp 1669390400
transform 1 0 104160 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_922
timestamp 1669390400
transform 1 0 104608 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_925
timestamp 1669390400
transform 1 0 104944 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_989
timestamp 1669390400
transform 1 0 112112 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_993
timestamp 1669390400
transform 1 0 112560 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_996
timestamp 1669390400
transform 1 0 112896 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_1030
timestamp 1669390400
transform 1 0 116704 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1038
timestamp 1669390400
transform 1 0 117600 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_1042
timestamp 1669390400
transform 1 0 118048 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1044
timestamp 1669390400
transform 1 0 118272 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_5
timestamp 1669390400
transform 1 0 1904 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_21
timestamp 1669390400
transform 1 0 3696 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_29
timestamp 1669390400
transform 1 0 4592 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_33
timestamp 1669390400
transform 1 0 5040 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1669390400
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1669390400
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1669390400
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1669390400
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1669390400
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1669390400
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_408
timestamp 1669390400
transform 1 0 47040 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_416
timestamp 1669390400
transform 1 0 47936 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_449
timestamp 1669390400
transform 1 0 51632 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_453
timestamp 1669390400
transform 1 0 52080 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_456
timestamp 1669390400
transform 1 0 52416 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_470
timestamp 1669390400
transform 1 0 53984 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_472
timestamp 1669390400
transform 1 0 54208 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_478
timestamp 1669390400
transform 1 0 54880 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_482
timestamp 1669390400
transform 1 0 55328 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_492
timestamp 1669390400
transform 1 0 56448 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_500
timestamp 1669390400
transform 1 0 57344 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_502
timestamp 1669390400
transform 1 0 57568 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_511
timestamp 1669390400
transform 1 0 58576 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_523
timestamp 1669390400
transform 1 0 59920 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_529
timestamp 1669390400
transform 1 0 60592 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1669390400
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_540
timestamp 1669390400
transform 1 0 61824 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_548
timestamp 1669390400
transform 1 0 62720 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_550
timestamp 1669390400
transform 1 0 62944 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_553
timestamp 1669390400
transform 1 0 63280 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_561
timestamp 1669390400
transform 1 0 64176 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_565
timestamp 1669390400
transform 1 0 64624 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_569
timestamp 1669390400
transform 1 0 65072 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_573
timestamp 1669390400
transform 1 0 65520 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_577
timestamp 1669390400
transform 1 0 65968 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_581
timestamp 1669390400
transform 1 0 66416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_585
timestamp 1669390400
transform 1 0 66864 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_587
timestamp 1669390400
transform 1 0 67088 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_590
timestamp 1669390400
transform 1 0 67424 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_594
timestamp 1669390400
transform 1 0 67872 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_598
timestamp 1669390400
transform 1 0 68320 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1669390400
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_605
timestamp 1669390400
transform 1 0 69104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_617
timestamp 1669390400
transform 1 0 70448 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_626
timestamp 1669390400
transform 1 0 71456 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_630
timestamp 1669390400
transform 1 0 71904 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_662
timestamp 1669390400
transform 1 0 75488 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_670
timestamp 1669390400
transform 1 0 76384 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_676
timestamp 1669390400
transform 1 0 77056 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_740
timestamp 1669390400
transform 1 0 84224 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_744
timestamp 1669390400
transform 1 0 84672 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_747
timestamp 1669390400
transform 1 0 85008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_811
timestamp 1669390400
transform 1 0 92176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_815
timestamp 1669390400
transform 1 0 92624 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_818
timestamp 1669390400
transform 1 0 92960 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_882
timestamp 1669390400
transform 1 0 100128 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_886
timestamp 1669390400
transform 1 0 100576 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_889
timestamp 1669390400
transform 1 0 100912 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_953
timestamp 1669390400
transform 1 0 108080 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_957
timestamp 1669390400
transform 1 0 108528 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_960
timestamp 1669390400
transform 1 0 108864 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_992
timestamp 1669390400
transform 1 0 112448 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1008
timestamp 1669390400
transform 1 0 114240 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1028
timestamp 1669390400
transform 1 0 116480 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1031
timestamp 1669390400
transform 1 0 116816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_1034
timestamp 1669390400
transform 1 0 117152 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_1042
timestamp 1669390400
transform 1 0 118048 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1044
timestamp 1669390400
transform 1 0 118272 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_19
timestamp 1669390400
transform 1 0 3472 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_51
timestamp 1669390400
transform 1 0 7056 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_67
timestamp 1669390400
transform 1 0 8848 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1669390400
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1669390400
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1669390400
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1669390400
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1669390400
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1669390400
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1669390400
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_421
timestamp 1669390400
transform 1 0 48496 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1669390400
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_435
timestamp 1669390400
transform 1 0 50064 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_439
timestamp 1669390400
transform 1 0 50512 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_469
timestamp 1669390400
transform 1 0 53872 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_481
timestamp 1669390400
transform 1 0 55216 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_493
timestamp 1669390400
transform 1 0 56560 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_505
timestamp 1669390400
transform 1 0 57904 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_517
timestamp 1669390400
transform 1 0 59248 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_527
timestamp 1669390400
transform 1 0 60368 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_529
timestamp 1669390400
transform 1 0 60592 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_536
timestamp 1669390400
transform 1 0 61376 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_540
timestamp 1669390400
transform 1 0 61824 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_544
timestamp 1669390400
transform 1 0 62272 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_560
timestamp 1669390400
transform 1 0 64064 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_564
timestamp 1669390400
transform 1 0 64512 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_570
timestamp 1669390400
transform 1 0 65184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_573
timestamp 1669390400
transform 1 0 65520 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_581
timestamp 1669390400
transform 1 0 66416 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_585
timestamp 1669390400
transform 1 0 66864 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_589
timestamp 1669390400
transform 1 0 67312 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_593
timestamp 1669390400
transform 1 0 67760 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_597
timestamp 1669390400
transform 1 0 68208 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_601
timestamp 1669390400
transform 1 0 68656 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_605
timestamp 1669390400
transform 1 0 69104 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_616
timestamp 1669390400
transform 1 0 70336 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_620
timestamp 1669390400
transform 1 0 70784 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_624
timestamp 1669390400
transform 1 0 71232 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_628
timestamp 1669390400
transform 1 0 71680 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_632
timestamp 1669390400
transform 1 0 72128 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_636
timestamp 1669390400
transform 1 0 72576 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1669390400
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_641
timestamp 1669390400
transform 1 0 73136 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_705
timestamp 1669390400
transform 1 0 80304 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_709
timestamp 1669390400
transform 1 0 80752 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_712
timestamp 1669390400
transform 1 0 81088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_776
timestamp 1669390400
transform 1 0 88256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_780
timestamp 1669390400
transform 1 0 88704 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_783
timestamp 1669390400
transform 1 0 89040 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_847
timestamp 1669390400
transform 1 0 96208 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_851
timestamp 1669390400
transform 1 0 96656 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_854
timestamp 1669390400
transform 1 0 96992 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_918
timestamp 1669390400
transform 1 0 104160 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_922
timestamp 1669390400
transform 1 0 104608 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_925
timestamp 1669390400
transform 1 0 104944 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_989
timestamp 1669390400
transform 1 0 112112 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_993
timestamp 1669390400
transform 1 0 112560 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_996
timestamp 1669390400
transform 1 0 112896 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_1028
timestamp 1669390400
transform 1 0 116480 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1044
timestamp 1669390400
transform 1 0 118272 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_19
timestamp 1669390400
transform 1 0 3472 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1669390400
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1669390400
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1669390400
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1669390400
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1669390400
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1669390400
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1669390400
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1669390400
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1669390400
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1669390400
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1669390400
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1669390400
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_392
timestamp 1669390400
transform 1 0 45248 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_400
timestamp 1669390400
transform 1 0 46144 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_402
timestamp 1669390400
transform 1 0 46368 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_405
timestamp 1669390400
transform 1 0 46704 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_409
timestamp 1669390400
transform 1 0 47152 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_413
timestamp 1669390400
transform 1 0 47600 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_417
timestamp 1669390400
transform 1 0 48048 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_421
timestamp 1669390400
transform 1 0 48496 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_425
timestamp 1669390400
transform 1 0 48944 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_441
timestamp 1669390400
transform 1 0 50736 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_445
timestamp 1669390400
transform 1 0 51184 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_448
timestamp 1669390400
transform 1 0 51520 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_452
timestamp 1669390400
transform 1 0 51968 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_456
timestamp 1669390400
transform 1 0 52416 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1669390400
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_463
timestamp 1669390400
transform 1 0 53200 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_472
timestamp 1669390400
transform 1 0 54208 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_476
timestamp 1669390400
transform 1 0 54656 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_488
timestamp 1669390400
transform 1 0 56000 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_499
timestamp 1669390400
transform 1 0 57232 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_506
timestamp 1669390400
transform 1 0 58016 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_514
timestamp 1669390400
transform 1 0 58912 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_526
timestamp 1669390400
transform 1 0 60256 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_530
timestamp 1669390400
transform 1 0 60704 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_537
timestamp 1669390400
transform 1 0 61488 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_539
timestamp 1669390400
transform 1 0 61712 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_542
timestamp 1669390400
transform 1 0 62048 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_546
timestamp 1669390400
transform 1 0 62496 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_550
timestamp 1669390400
transform 1 0 62944 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_552
timestamp 1669390400
transform 1 0 63168 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_584
timestamp 1669390400
transform 1 0 66752 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_588
timestamp 1669390400
transform 1 0 67200 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_592
timestamp 1669390400
transform 1 0 67648 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_594
timestamp 1669390400
transform 1 0 67872 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1669390400
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_605
timestamp 1669390400
transform 1 0 69104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_615
timestamp 1669390400
transform 1 0 70224 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_619
timestamp 1669390400
transform 1 0 70672 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_623
timestamp 1669390400
transform 1 0 71120 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_627
timestamp 1669390400
transform 1 0 71568 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_631
timestamp 1669390400
transform 1 0 72016 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_639
timestamp 1669390400
transform 1 0 72912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_642
timestamp 1669390400
transform 1 0 73248 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_676
timestamp 1669390400
transform 1 0 77056 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_740
timestamp 1669390400
transform 1 0 84224 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_744
timestamp 1669390400
transform 1 0 84672 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_747
timestamp 1669390400
transform 1 0 85008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_811
timestamp 1669390400
transform 1 0 92176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_815
timestamp 1669390400
transform 1 0 92624 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_818
timestamp 1669390400
transform 1 0 92960 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_882
timestamp 1669390400
transform 1 0 100128 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_886
timestamp 1669390400
transform 1 0 100576 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_889
timestamp 1669390400
transform 1 0 100912 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_953
timestamp 1669390400
transform 1 0 108080 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_957
timestamp 1669390400
transform 1 0 108528 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_960
timestamp 1669390400
transform 1 0 108864 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_992
timestamp 1669390400
transform 1 0 112448 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1008
timestamp 1669390400
transform 1 0 114240 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1012
timestamp 1669390400
transform 1 0 114688 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_1019
timestamp 1669390400
transform 1 0 115472 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1023
timestamp 1669390400
transform 1 0 115920 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_1027
timestamp 1669390400
transform 1 0 116368 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_1031
timestamp 1669390400
transform 1 0 116816 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1039
timestamp 1669390400
transform 1 0 117712 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_1043
timestamp 1669390400
transform 1 0 118160 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_5
timestamp 1669390400
transform 1 0 1904 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_69
timestamp 1669390400
transform 1 0 9072 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1669390400
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1669390400
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1669390400
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1669390400
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1669390400
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1669390400
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1669390400
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1669390400
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1669390400
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1669390400
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1669390400
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_357
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_389
timestamp 1669390400
transform 1 0 44912 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_393
timestamp 1669390400
transform 1 0 45360 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_409
timestamp 1669390400
transform 1 0 47152 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1669390400
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_428
timestamp 1669390400
transform 1 0 49280 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_441
timestamp 1669390400
transform 1 0 50736 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_445
timestamp 1669390400
transform 1 0 51184 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_449
timestamp 1669390400
transform 1 0 51632 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_455
timestamp 1669390400
transform 1 0 52304 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_459
timestamp 1669390400
transform 1 0 52752 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_463
timestamp 1669390400
transform 1 0 53200 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_467
timestamp 1669390400
transform 1 0 53648 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_475
timestamp 1669390400
transform 1 0 54544 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_485
timestamp 1669390400
transform 1 0 55664 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_493
timestamp 1669390400
transform 1 0 56560 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_499
timestamp 1669390400
transform 1 0 57232 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_505
timestamp 1669390400
transform 1 0 57904 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_513
timestamp 1669390400
transform 1 0 58800 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_524
timestamp 1669390400
transform 1 0 60032 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_528
timestamp 1669390400
transform 1 0 60480 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_532
timestamp 1669390400
transform 1 0 60928 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_534
timestamp 1669390400
transform 1 0 61152 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_543
timestamp 1669390400
transform 1 0 62160 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_547
timestamp 1669390400
transform 1 0 62608 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_561
timestamp 1669390400
transform 1 0 64176 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_565
timestamp 1669390400
transform 1 0 64624 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1669390400
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_570
timestamp 1669390400
transform 1 0 65184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_577
timestamp 1669390400
transform 1 0 65968 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_581
timestamp 1669390400
transform 1 0 66416 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_585
timestamp 1669390400
transform 1 0 66864 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_597
timestamp 1669390400
transform 1 0 68208 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_603
timestamp 1669390400
transform 1 0 68880 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_618
timestamp 1669390400
transform 1 0 70560 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_624
timestamp 1669390400
transform 1 0 71232 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_626
timestamp 1669390400
transform 1 0 71456 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_635
timestamp 1669390400
transform 1 0 72464 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_641
timestamp 1669390400
transform 1 0 73136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_648
timestamp 1669390400
transform 1 0 73920 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_652
timestamp 1669390400
transform 1 0 74368 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_684
timestamp 1669390400
transform 1 0 77952 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_700
timestamp 1669390400
transform 1 0 79744 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_708
timestamp 1669390400
transform 1 0 80640 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_712
timestamp 1669390400
transform 1 0 81088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_776
timestamp 1669390400
transform 1 0 88256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_780
timestamp 1669390400
transform 1 0 88704 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_783
timestamp 1669390400
transform 1 0 89040 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_847
timestamp 1669390400
transform 1 0 96208 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_851
timestamp 1669390400
transform 1 0 96656 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_854
timestamp 1669390400
transform 1 0 96992 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_918
timestamp 1669390400
transform 1 0 104160 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_922
timestamp 1669390400
transform 1 0 104608 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_925
timestamp 1669390400
transform 1 0 104944 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_989
timestamp 1669390400
transform 1 0 112112 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_993
timestamp 1669390400
transform 1 0 112560 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_996
timestamp 1669390400
transform 1 0 112896 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1012
timestamp 1669390400
transform 1 0 114688 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_1029
timestamp 1669390400
transform 1 0 116592 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_1033
timestamp 1669390400
transform 1 0 117040 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1041
timestamp 1669390400
transform 1 0 117936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_17
timestamp 1669390400
transform 1 0 3248 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_21
timestamp 1669390400
transform 1 0 3696 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_29
timestamp 1669390400
transform 1 0 4592 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_33
timestamp 1669390400
transform 1 0 5040 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1669390400
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1669390400
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1669390400
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1669390400
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1669390400
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1669390400
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1669390400
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1669390400
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1669390400
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1669390400
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1669390400
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1669390400
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1669390400
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1669390400
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1669390400
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_392
timestamp 1669390400
transform 1 0 45248 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_422
timestamp 1669390400
transform 1 0 48608 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_426
timestamp 1669390400
transform 1 0 49056 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_430
timestamp 1669390400
transform 1 0 49504 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_438
timestamp 1669390400
transform 1 0 50400 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_440
timestamp 1669390400
transform 1 0 50624 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_443
timestamp 1669390400
transform 1 0 50960 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_447
timestamp 1669390400
transform 1 0 51408 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_451
timestamp 1669390400
transform 1 0 51856 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_453
timestamp 1669390400
transform 1 0 52080 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_456
timestamp 1669390400
transform 1 0 52416 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1669390400
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_463
timestamp 1669390400
transform 1 0 53200 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_467
timestamp 1669390400
transform 1 0 53648 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_475
timestamp 1669390400
transform 1 0 54544 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_481
timestamp 1669390400
transform 1 0 55216 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_485
timestamp 1669390400
transform 1 0 55664 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_489
timestamp 1669390400
transform 1 0 56112 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_493
timestamp 1669390400
transform 1 0 56560 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_497
timestamp 1669390400
transform 1 0 57008 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_503
timestamp 1669390400
transform 1 0 57680 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_507
timestamp 1669390400
transform 1 0 58128 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_511
timestamp 1669390400
transform 1 0 58576 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_515
timestamp 1669390400
transform 1 0 59024 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_519
timestamp 1669390400
transform 1 0 59472 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_523
timestamp 1669390400
transform 1 0 59920 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1669390400
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_585
timestamp 1669390400
transform 1 0 66864 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_596
timestamp 1669390400
transform 1 0 68096 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_600
timestamp 1669390400
transform 1 0 68544 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1669390400
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_605
timestamp 1669390400
transform 1 0 69104 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_607
timestamp 1669390400
transform 1 0 69328 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_616
timestamp 1669390400
transform 1 0 70336 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_618
timestamp 1669390400
transform 1 0 70560 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_623
timestamp 1669390400
transform 1 0 71120 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_625
timestamp 1669390400
transform 1 0 71344 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_655
timestamp 1669390400
transform 1 0 74704 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_659
timestamp 1669390400
transform 1 0 75152 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_667
timestamp 1669390400
transform 1 0 76048 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_671
timestamp 1669390400
transform 1 0 76496 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1669390400
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_676
timestamp 1669390400
transform 1 0 77056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_727
timestamp 1669390400
transform 1 0 82768 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_731
timestamp 1669390400
transform 1 0 83216 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_739
timestamp 1669390400
transform 1 0 84112 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_743
timestamp 1669390400
transform 1 0 84560 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_747
timestamp 1669390400
transform 1 0 85008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_811
timestamp 1669390400
transform 1 0 92176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_815
timestamp 1669390400
transform 1 0 92624 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_818
timestamp 1669390400
transform 1 0 92960 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_882
timestamp 1669390400
transform 1 0 100128 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_886
timestamp 1669390400
transform 1 0 100576 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_889
timestamp 1669390400
transform 1 0 100912 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_953
timestamp 1669390400
transform 1 0 108080 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_957
timestamp 1669390400
transform 1 0 108528 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_960
timestamp 1669390400
transform 1 0 108864 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_992
timestamp 1669390400
transform 1 0 112448 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1008
timestamp 1669390400
transform 1 0 114240 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1028
timestamp 1669390400
transform 1 0 116480 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1031
timestamp 1669390400
transform 1 0 116816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_1034
timestamp 1669390400
transform 1 0 117152 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_1042
timestamp 1669390400
transform 1 0 118048 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1044
timestamp 1669390400
transform 1 0 118272 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_5
timestamp 1669390400
transform 1 0 1904 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_69
timestamp 1669390400
transform 1 0 9072 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1669390400
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1669390400
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1669390400
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1669390400
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1669390400
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1669390400
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1669390400
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1669390400
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1669390400
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1669390400
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1669390400
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_357
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_389
timestamp 1669390400
transform 1 0 44912 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_399
timestamp 1669390400
transform 1 0 46032 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_415
timestamp 1669390400
transform 1 0 47824 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1669390400
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1669390400
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_428
timestamp 1669390400
transform 1 0 49280 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_432
timestamp 1669390400
transform 1 0 49728 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_442
timestamp 1669390400
transform 1 0 50848 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_446
timestamp 1669390400
transform 1 0 51296 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_454
timestamp 1669390400
transform 1 0 52192 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_458
timestamp 1669390400
transform 1 0 52640 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_461
timestamp 1669390400
transform 1 0 52976 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_465
timestamp 1669390400
transform 1 0 53424 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_471
timestamp 1669390400
transform 1 0 54096 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_487
timestamp 1669390400
transform 1 0 55888 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_489
timestamp 1669390400
transform 1 0 56112 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_492
timestamp 1669390400
transform 1 0 56448 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1669390400
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_499
timestamp 1669390400
transform 1 0 57232 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_512
timestamp 1669390400
transform 1 0 58688 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_516
timestamp 1669390400
transform 1 0 59136 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_549
timestamp 1669390400
transform 1 0 62832 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_553
timestamp 1669390400
transform 1 0 63280 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_563
timestamp 1669390400
transform 1 0 64400 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1669390400
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_570
timestamp 1669390400
transform 1 0 65184 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_577
timestamp 1669390400
transform 1 0 65968 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_581
timestamp 1669390400
transform 1 0 66416 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_611
timestamp 1669390400
transform 1 0 69776 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_615
timestamp 1669390400
transform 1 0 70224 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_619
timestamp 1669390400
transform 1 0 70672 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_623
timestamp 1669390400
transform 1 0 71120 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_627
timestamp 1669390400
transform 1 0 71568 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_636
timestamp 1669390400
transform 1 0 72576 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1669390400
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_641
timestamp 1669390400
transform 1 0 73136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_648
timestamp 1669390400
transform 1 0 73920 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_652
timestamp 1669390400
transform 1 0 74368 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_656
timestamp 1669390400
transform 1 0 74816 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_688
timestamp 1669390400
transform 1 0 78400 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_704
timestamp 1669390400
transform 1 0 80192 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_708
timestamp 1669390400
transform 1 0 80640 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_712
timestamp 1669390400
transform 1 0 81088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_776
timestamp 1669390400
transform 1 0 88256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_780
timestamp 1669390400
transform 1 0 88704 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_783
timestamp 1669390400
transform 1 0 89040 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_847
timestamp 1669390400
transform 1 0 96208 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_851
timestamp 1669390400
transform 1 0 96656 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_854
timestamp 1669390400
transform 1 0 96992 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_918
timestamp 1669390400
transform 1 0 104160 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_922
timestamp 1669390400
transform 1 0 104608 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_925
timestamp 1669390400
transform 1 0 104944 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_989
timestamp 1669390400
transform 1 0 112112 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_993
timestamp 1669390400
transform 1 0 112560 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_996
timestamp 1669390400
transform 1 0 112896 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_1028
timestamp 1669390400
transform 1 0 116480 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1044
timestamp 1669390400
transform 1 0 118272 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_19
timestamp 1669390400
transform 1 0 3472 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1669390400
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1669390400
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1669390400
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1669390400
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1669390400
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1669390400
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1669390400
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1669390400
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1669390400
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1669390400
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1669390400
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1669390400
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1669390400
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1669390400
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1669390400
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_392
timestamp 1669390400
transform 1 0 45248 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_408
timestamp 1669390400
transform 1 0 47040 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_410
timestamp 1669390400
transform 1 0 47264 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_419
timestamp 1669390400
transform 1 0 48272 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_450
timestamp 1669390400
transform 1 0 51744 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_454
timestamp 1669390400
transform 1 0 52192 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_458
timestamp 1669390400
transform 1 0 52640 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1669390400
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_463
timestamp 1669390400
transform 1 0 53200 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_495
timestamp 1669390400
transform 1 0 56784 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_499
timestamp 1669390400
transform 1 0 57232 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_502
timestamp 1669390400
transform 1 0 57568 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_518
timestamp 1669390400
transform 1 0 59360 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_522
timestamp 1669390400
transform 1 0 59808 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_530
timestamp 1669390400
transform 1 0 60704 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_538
timestamp 1669390400
transform 1 0 61600 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_545
timestamp 1669390400
transform 1 0 62384 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_547
timestamp 1669390400
transform 1 0 62608 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_554
timestamp 1669390400
transform 1 0 63392 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_593
timestamp 1669390400
transform 1 0 67760 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_597
timestamp 1669390400
transform 1 0 68208 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_601
timestamp 1669390400
transform 1 0 68656 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_605
timestamp 1669390400
transform 1 0 69104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_612
timestamp 1669390400
transform 1 0 69888 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_616
timestamp 1669390400
transform 1 0 70336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_620
timestamp 1669390400
transform 1 0 70784 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_624
timestamp 1669390400
transform 1 0 71232 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_655
timestamp 1669390400
transform 1 0 74704 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_659
timestamp 1669390400
transform 1 0 75152 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_667
timestamp 1669390400
transform 1 0 76048 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_671
timestamp 1669390400
transform 1 0 76496 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1669390400
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_676
timestamp 1669390400
transform 1 0 77056 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_740
timestamp 1669390400
transform 1 0 84224 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_744
timestamp 1669390400
transform 1 0 84672 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_747
timestamp 1669390400
transform 1 0 85008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_811
timestamp 1669390400
transform 1 0 92176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_815
timestamp 1669390400
transform 1 0 92624 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_818
timestamp 1669390400
transform 1 0 92960 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_882
timestamp 1669390400
transform 1 0 100128 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_886
timestamp 1669390400
transform 1 0 100576 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_889
timestamp 1669390400
transform 1 0 100912 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_953
timestamp 1669390400
transform 1 0 108080 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_957
timestamp 1669390400
transform 1 0 108528 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_960
timestamp 1669390400
transform 1 0 108864 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_992
timestamp 1669390400
transform 1 0 112448 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1008
timestamp 1669390400
transform 1 0 114240 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1028
timestamp 1669390400
transform 1 0 116480 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1031
timestamp 1669390400
transform 1 0 116816 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_1034
timestamp 1669390400
transform 1 0 117152 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_1042
timestamp 1669390400
transform 1 0 118048 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1044
timestamp 1669390400
transform 1 0 118272 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_19
timestamp 1669390400
transform 1 0 3472 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_51
timestamp 1669390400
transform 1 0 7056 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_67
timestamp 1669390400
transform 1 0 8848 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1669390400
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1669390400
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1669390400
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1669390400
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1669390400
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1669390400
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1669390400
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1669390400
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1669390400
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1669390400
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1669390400
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_357
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_389
timestamp 1669390400
transform 1 0 44912 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_393
timestamp 1669390400
transform 1 0 45360 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_395
timestamp 1669390400
transform 1 0 45584 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1669390400
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_428
timestamp 1669390400
transform 1 0 49280 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_435
timestamp 1669390400
transform 1 0 50064 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_443
timestamp 1669390400
transform 1 0 50960 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_447
timestamp 1669390400
transform 1 0 51408 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_463
timestamp 1669390400
transform 1 0 53200 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_467
timestamp 1669390400
transform 1 0 53648 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_475
timestamp 1669390400
transform 1 0 54544 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_489
timestamp 1669390400
transform 1 0 56112 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_493
timestamp 1669390400
transform 1 0 56560 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1669390400
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_499
timestamp 1669390400
transform 1 0 57232 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_501
timestamp 1669390400
transform 1 0 57456 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_504
timestamp 1669390400
transform 1 0 57792 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_512
timestamp 1669390400
transform 1 0 58688 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_543
timestamp 1669390400
transform 1 0 62160 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_553
timestamp 1669390400
transform 1 0 63280 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_563
timestamp 1669390400
transform 1 0 64400 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1669390400
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_570
timestamp 1669390400
transform 1 0 65184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_576
timestamp 1669390400
transform 1 0 65856 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_580
timestamp 1669390400
transform 1 0 66304 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_584
timestamp 1669390400
transform 1 0 66752 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_594
timestamp 1669390400
transform 1 0 67872 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_598
timestamp 1669390400
transform 1 0 68320 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_602
timestamp 1669390400
transform 1 0 68768 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_606
timestamp 1669390400
transform 1 0 69216 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_610
timestamp 1669390400
transform 1 0 69664 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_614
timestamp 1669390400
transform 1 0 70112 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_621
timestamp 1669390400
transform 1 0 70896 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_625
timestamp 1669390400
transform 1 0 71344 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_633
timestamp 1669390400
transform 1 0 72240 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_637
timestamp 1669390400
transform 1 0 72688 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_641
timestamp 1669390400
transform 1 0 73136 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_705
timestamp 1669390400
transform 1 0 80304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_709
timestamp 1669390400
transform 1 0 80752 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_712
timestamp 1669390400
transform 1 0 81088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_776
timestamp 1669390400
transform 1 0 88256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_780
timestamp 1669390400
transform 1 0 88704 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_783
timestamp 1669390400
transform 1 0 89040 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_847
timestamp 1669390400
transform 1 0 96208 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_851
timestamp 1669390400
transform 1 0 96656 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_854
timestamp 1669390400
transform 1 0 96992 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_918
timestamp 1669390400
transform 1 0 104160 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_922
timestamp 1669390400
transform 1 0 104608 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_925
timestamp 1669390400
transform 1 0 104944 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_989
timestamp 1669390400
transform 1 0 112112 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_993
timestamp 1669390400
transform 1 0 112560 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_996
timestamp 1669390400
transform 1 0 112896 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_1028
timestamp 1669390400
transform 1 0 116480 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1044
timestamp 1669390400
transform 1 0 118272 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_5
timestamp 1669390400
transform 1 0 1904 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_21
timestamp 1669390400
transform 1 0 3696 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_29
timestamp 1669390400
transform 1 0 4592 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_33
timestamp 1669390400
transform 1 0 5040 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1669390400
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1669390400
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1669390400
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1669390400
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1669390400
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1669390400
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1669390400
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1669390400
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1669390400
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1669390400
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1669390400
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1669390400
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1669390400
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_385
timestamp 1669390400
transform 1 0 44464 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1669390400
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_392
timestamp 1669390400
transform 1 0 45248 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_408
timestamp 1669390400
transform 1 0 47040 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_412
timestamp 1669390400
transform 1 0 47488 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_422
timestamp 1669390400
transform 1 0 48608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_426
timestamp 1669390400
transform 1 0 49056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_429
timestamp 1669390400
transform 1 0 49392 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_433
timestamp 1669390400
transform 1 0 49840 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_437
timestamp 1669390400
transform 1 0 50288 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_441
timestamp 1669390400
transform 1 0 50736 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_457
timestamp 1669390400
transform 1 0 52528 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_463
timestamp 1669390400
transform 1 0 53200 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_471
timestamp 1669390400
transform 1 0 54096 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_474
timestamp 1669390400
transform 1 0 54432 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_476
timestamp 1669390400
transform 1 0 54656 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_479
timestamp 1669390400
transform 1 0 54992 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_483
timestamp 1669390400
transform 1 0 55440 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_487
timestamp 1669390400
transform 1 0 55888 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_521
timestamp 1669390400
transform 1 0 59696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_527
timestamp 1669390400
transform 1 0 60368 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1669390400
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_542
timestamp 1669390400
transform 1 0 62048 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_545
timestamp 1669390400
transform 1 0 62384 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_549
timestamp 1669390400
transform 1 0 62832 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_565
timestamp 1669390400
transform 1 0 64624 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_569
timestamp 1669390400
transform 1 0 65072 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_574
timestamp 1669390400
transform 1 0 65632 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_576
timestamp 1669390400
transform 1 0 65856 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_585
timestamp 1669390400
transform 1 0 66864 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_589
timestamp 1669390400
transform 1 0 67312 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_597
timestamp 1669390400
transform 1 0 68208 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_601
timestamp 1669390400
transform 1 0 68656 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_605
timestamp 1669390400
transform 1 0 69104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_614
timestamp 1669390400
transform 1 0 70112 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_622
timestamp 1669390400
transform 1 0 71008 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_626
timestamp 1669390400
transform 1 0 71456 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_630
timestamp 1669390400
transform 1 0 71904 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_634
timestamp 1669390400
transform 1 0 72352 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_666
timestamp 1669390400
transform 1 0 75936 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_676
timestamp 1669390400
transform 1 0 77056 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_740
timestamp 1669390400
transform 1 0 84224 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_744
timestamp 1669390400
transform 1 0 84672 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_747
timestamp 1669390400
transform 1 0 85008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_811
timestamp 1669390400
transform 1 0 92176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_815
timestamp 1669390400
transform 1 0 92624 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_818
timestamp 1669390400
transform 1 0 92960 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_882
timestamp 1669390400
transform 1 0 100128 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_886
timestamp 1669390400
transform 1 0 100576 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_889
timestamp 1669390400
transform 1 0 100912 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_953
timestamp 1669390400
transform 1 0 108080 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_957
timestamp 1669390400
transform 1 0 108528 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_960
timestamp 1669390400
transform 1 0 108864 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_992
timestamp 1669390400
transform 1 0 112448 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1008
timestamp 1669390400
transform 1 0 114240 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1028
timestamp 1669390400
transform 1 0 116480 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1031
timestamp 1669390400
transform 1 0 116816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_1034
timestamp 1669390400
transform 1 0 117152 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_1042
timestamp 1669390400
transform 1 0 118048 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1044
timestamp 1669390400
transform 1 0 118272 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_5
timestamp 1669390400
transform 1 0 1904 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_69
timestamp 1669390400
transform 1 0 9072 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1669390400
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1669390400
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1669390400
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1669390400
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1669390400
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1669390400
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1669390400
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1669390400
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1669390400
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1669390400
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1669390400
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_357
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_373
timestamp 1669390400
transform 1 0 43120 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_381
timestamp 1669390400
transform 1 0 44016 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_414
timestamp 1669390400
transform 1 0 47712 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_418
timestamp 1669390400
transform 1 0 48160 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_424
timestamp 1669390400
transform 1 0 48832 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_428
timestamp 1669390400
transform 1 0 49280 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_431
timestamp 1669390400
transform 1 0 49616 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_435
timestamp 1669390400
transform 1 0 50064 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_451
timestamp 1669390400
transform 1 0 51856 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_459
timestamp 1669390400
transform 1 0 52752 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_465
timestamp 1669390400
transform 1 0 53424 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_469
timestamp 1669390400
transform 1 0 53872 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_473
timestamp 1669390400
transform 1 0 54320 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_477
timestamp 1669390400
transform 1 0 54768 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_481
timestamp 1669390400
transform 1 0 55216 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_491
timestamp 1669390400
transform 1 0 56336 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_495
timestamp 1669390400
transform 1 0 56784 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_499
timestamp 1669390400
transform 1 0 57232 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_502
timestamp 1669390400
transform 1 0 57568 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_508
timestamp 1669390400
transform 1 0 58240 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_512
timestamp 1669390400
transform 1 0 58688 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_520
timestamp 1669390400
transform 1 0 59584 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_523
timestamp 1669390400
transform 1 0 59920 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_531
timestamp 1669390400
transform 1 0 60816 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_534
timestamp 1669390400
transform 1 0 61152 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_538
timestamp 1669390400
transform 1 0 61600 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_556
timestamp 1669390400
transform 1 0 63616 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_560
timestamp 1669390400
transform 1 0 64064 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_564
timestamp 1669390400
transform 1 0 64512 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1669390400
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_570
timestamp 1669390400
transform 1 0 65184 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_572
timestamp 1669390400
transform 1 0 65408 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_602
timestamp 1669390400
transform 1 0 68768 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_633
timestamp 1669390400
transform 1 0 72240 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_637
timestamp 1669390400
transform 1 0 72688 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_641
timestamp 1669390400
transform 1 0 73136 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_649
timestamp 1669390400
transform 1 0 74032 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_652
timestamp 1669390400
transform 1 0 74368 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_656
timestamp 1669390400
transform 1 0 74816 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_660
timestamp 1669390400
transform 1 0 75264 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_676
timestamp 1669390400
transform 1 0 77056 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_678
timestamp 1669390400
transform 1 0 77280 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_681
timestamp 1669390400
transform 1 0 77616 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_697
timestamp 1669390400
transform 1 0 79408 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_705
timestamp 1669390400
transform 1 0 80304 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_709
timestamp 1669390400
transform 1 0 80752 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_712
timestamp 1669390400
transform 1 0 81088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_776
timestamp 1669390400
transform 1 0 88256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_780
timestamp 1669390400
transform 1 0 88704 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_783
timestamp 1669390400
transform 1 0 89040 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_847
timestamp 1669390400
transform 1 0 96208 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_851
timestamp 1669390400
transform 1 0 96656 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_854
timestamp 1669390400
transform 1 0 96992 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_918
timestamp 1669390400
transform 1 0 104160 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_922
timestamp 1669390400
transform 1 0 104608 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_925
timestamp 1669390400
transform 1 0 104944 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_989
timestamp 1669390400
transform 1 0 112112 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_993
timestamp 1669390400
transform 1 0 112560 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_996
timestamp 1669390400
transform 1 0 112896 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1004
timestamp 1669390400
transform 1 0 113792 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_1007
timestamp 1669390400
transform 1 0 114128 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_1038
timestamp 1669390400
transform 1 0 117600 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_1042
timestamp 1669390400
transform 1 0 118048 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1044
timestamp 1669390400
transform 1 0 118272 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_19
timestamp 1669390400
transform 1 0 3472 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1669390400
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1669390400
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1669390400
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1669390400
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1669390400
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1669390400
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1669390400
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1669390400
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1669390400
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1669390400
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1669390400
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1669390400
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1669390400
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1669390400
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1669390400
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_392
timestamp 1669390400
transform 1 0 45248 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_399
timestamp 1669390400
transform 1 0 46032 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_407
timestamp 1669390400
transform 1 0 46928 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_438
timestamp 1669390400
transform 1 0 50400 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_442
timestamp 1669390400
transform 1 0 50848 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_452
timestamp 1669390400
transform 1 0 51968 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1669390400
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_463
timestamp 1669390400
transform 1 0 53200 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_465
timestamp 1669390400
transform 1 0 53424 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_472
timestamp 1669390400
transform 1 0 54208 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_488
timestamp 1669390400
transform 1 0 56000 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_504
timestamp 1669390400
transform 1 0 57792 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_512
timestamp 1669390400
transform 1 0 58688 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_516
timestamp 1669390400
transform 1 0 59136 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_520
timestamp 1669390400
transform 1 0 59584 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_528
timestamp 1669390400
transform 1 0 60480 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1669390400
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_541
timestamp 1669390400
transform 1 0 61936 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_545
timestamp 1669390400
transform 1 0 62384 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_578
timestamp 1669390400
transform 1 0 66080 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_582
timestamp 1669390400
transform 1 0 66528 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_586
timestamp 1669390400
transform 1 0 66976 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_588
timestamp 1669390400
transform 1 0 67200 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_591
timestamp 1669390400
transform 1 0 67536 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_599
timestamp 1669390400
transform 1 0 68432 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_605
timestamp 1669390400
transform 1 0 69104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_608
timestamp 1669390400
transform 1 0 69440 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_616
timestamp 1669390400
transform 1 0 70336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_620
timestamp 1669390400
transform 1 0 70784 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_622
timestamp 1669390400
transform 1 0 71008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_652
timestamp 1669390400
transform 1 0 74368 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_669
timestamp 1669390400
transform 1 0 76272 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1669390400
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_676
timestamp 1669390400
transform 1 0 77056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_679
timestamp 1669390400
transform 1 0 77392 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_696
timestamp 1669390400
transform 1 0 79296 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_700
timestamp 1669390400
transform 1 0 79744 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_716
timestamp 1669390400
transform 1 0 81536 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_719
timestamp 1669390400
transform 1 0 81872 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_735
timestamp 1669390400
transform 1 0 83664 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_743
timestamp 1669390400
transform 1 0 84560 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_747
timestamp 1669390400
transform 1 0 85008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_811
timestamp 1669390400
transform 1 0 92176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_815
timestamp 1669390400
transform 1 0 92624 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_818
timestamp 1669390400
transform 1 0 92960 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_882
timestamp 1669390400
transform 1 0 100128 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_886
timestamp 1669390400
transform 1 0 100576 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_889
timestamp 1669390400
transform 1 0 100912 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_953
timestamp 1669390400
transform 1 0 108080 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_957
timestamp 1669390400
transform 1 0 108528 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_960
timestamp 1669390400
transform 1 0 108864 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_992
timestamp 1669390400
transform 1 0 112448 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1000
timestamp 1669390400
transform 1 0 113344 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_1003
timestamp 1669390400
transform 1 0 113680 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_1011
timestamp 1669390400
transform 1 0 114576 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1028
timestamp 1669390400
transform 1 0 116480 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1031
timestamp 1669390400
transform 1 0 116816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_1038
timestamp 1669390400
transform 1 0 117600 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_1042
timestamp 1669390400
transform 1 0 118048 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1044
timestamp 1669390400
transform 1 0 118272 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_66
timestamp 1669390400
transform 1 0 8736 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1669390400
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1669390400
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1669390400
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1669390400
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1669390400
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1669390400
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1669390400
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1669390400
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1669390400
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1669390400
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1669390400
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1669390400
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_357
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_389
timestamp 1669390400
transform 1 0 44912 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_405
timestamp 1669390400
transform 1 0 46704 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_413
timestamp 1669390400
transform 1 0 47600 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_417
timestamp 1669390400
transform 1 0 48048 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_424
timestamp 1669390400
transform 1 0 48832 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_428
timestamp 1669390400
transform 1 0 49280 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_444
timestamp 1669390400
transform 1 0 51072 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_448
timestamp 1669390400
transform 1 0 51520 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_487
timestamp 1669390400
transform 1 0 55888 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_494
timestamp 1669390400
transform 1 0 56672 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1669390400
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_499
timestamp 1669390400
transform 1 0 57232 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_531
timestamp 1669390400
transform 1 0 60816 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_562
timestamp 1669390400
transform 1 0 64288 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_566
timestamp 1669390400
transform 1 0 64736 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_570
timestamp 1669390400
transform 1 0 65184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_573
timestamp 1669390400
transform 1 0 65520 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_605
timestamp 1669390400
transform 1 0 69104 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_613
timestamp 1669390400
transform 1 0 70000 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_617
timestamp 1669390400
transform 1 0 70448 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_621
timestamp 1669390400
transform 1 0 70896 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1669390400
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_641
timestamp 1669390400
transform 1 0 73136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_644
timestamp 1669390400
transform 1 0 73472 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_648
timestamp 1669390400
transform 1 0 73920 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_678
timestamp 1669390400
transform 1 0 77280 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_709
timestamp 1669390400
transform 1 0 80752 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_712
timestamp 1669390400
transform 1 0 81088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_715
timestamp 1669390400
transform 1 0 81424 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_725
timestamp 1669390400
transform 1 0 82544 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_757
timestamp 1669390400
transform 1 0 86128 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_773
timestamp 1669390400
transform 1 0 87920 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_783
timestamp 1669390400
transform 1 0 89040 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_847
timestamp 1669390400
transform 1 0 96208 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_851
timestamp 1669390400
transform 1 0 96656 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_854
timestamp 1669390400
transform 1 0 96992 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_918
timestamp 1669390400
transform 1 0 104160 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_922
timestamp 1669390400
transform 1 0 104608 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_925
timestamp 1669390400
transform 1 0 104944 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_989
timestamp 1669390400
transform 1 0 112112 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_993
timestamp 1669390400
transform 1 0 112560 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_996
timestamp 1669390400
transform 1 0 112896 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1004
timestamp 1669390400
transform 1 0 113792 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_1007
timestamp 1669390400
transform 1 0 114128 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1011
timestamp 1669390400
transform 1 0 114576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1044
timestamp 1669390400
transform 1 0 118272 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1669390400
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1669390400
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1669390400
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1669390400
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1669390400
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1669390400
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1669390400
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1669390400
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1669390400
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1669390400
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1669390400
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1669390400
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1669390400
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1669390400
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1669390400
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1669390400
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_392
timestamp 1669390400
transform 1 0 45248 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_424
timestamp 1669390400
transform 1 0 48832 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_426
timestamp 1669390400
transform 1 0 49056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_429
timestamp 1669390400
transform 1 0 49392 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_433
timestamp 1669390400
transform 1 0 49840 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_449
timestamp 1669390400
transform 1 0 51632 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_457
timestamp 1669390400
transform 1 0 52528 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_463
timestamp 1669390400
transform 1 0 53200 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_471
timestamp 1669390400
transform 1 0 54096 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_487
timestamp 1669390400
transform 1 0 55888 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_502
timestamp 1669390400
transform 1 0 57568 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_506
timestamp 1669390400
transform 1 0 58016 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_522
timestamp 1669390400
transform 1 0 59808 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_526
timestamp 1669390400
transform 1 0 60256 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_528
timestamp 1669390400
transform 1 0 60480 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1669390400
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_550
timestamp 1669390400
transform 1 0 62944 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_558
timestamp 1669390400
transform 1 0 63840 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_562
timestamp 1669390400
transform 1 0 64288 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_566
timestamp 1669390400
transform 1 0 64736 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_598
timestamp 1669390400
transform 1 0 68320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1669390400
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_605
timestamp 1669390400
transform 1 0 69104 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_621
timestamp 1669390400
transform 1 0 70896 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_625
timestamp 1669390400
transform 1 0 71344 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_633
timestamp 1669390400
transform 1 0 72240 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_649
timestamp 1669390400
transform 1 0 74032 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_653
timestamp 1669390400
transform 1 0 74480 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_660
timestamp 1669390400
transform 1 0 75264 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_668
timestamp 1669390400
transform 1 0 76160 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_672
timestamp 1669390400
transform 1 0 76608 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_676
timestamp 1669390400
transform 1 0 77056 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_684
timestamp 1669390400
transform 1 0 77952 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_688
timestamp 1669390400
transform 1 0 78400 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_720
timestamp 1669390400
transform 1 0 81984 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_736
timestamp 1669390400
transform 1 0 83776 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_744
timestamp 1669390400
transform 1 0 84672 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_747
timestamp 1669390400
transform 1 0 85008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_811
timestamp 1669390400
transform 1 0 92176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_815
timestamp 1669390400
transform 1 0 92624 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_818
timestamp 1669390400
transform 1 0 92960 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_882
timestamp 1669390400
transform 1 0 100128 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_886
timestamp 1669390400
transform 1 0 100576 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_889
timestamp 1669390400
transform 1 0 100912 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_953
timestamp 1669390400
transform 1 0 108080 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_957
timestamp 1669390400
transform 1 0 108528 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_960
timestamp 1669390400
transform 1 0 108864 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_992
timestamp 1669390400
transform 1 0 112448 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1008
timestamp 1669390400
transform 1 0 114240 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1012
timestamp 1669390400
transform 1 0 114688 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_1027
timestamp 1669390400
transform 1 0 116368 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1031
timestamp 1669390400
transform 1 0 116816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1038
timestamp 1669390400
transform 1 0 117600 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_1042
timestamp 1669390400
transform 1 0 118048 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1044
timestamp 1669390400
transform 1 0 118272 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_17
timestamp 1669390400
transform 1 0 3248 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_21
timestamp 1669390400
transform 1 0 3696 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_53
timestamp 1669390400
transform 1 0 7280 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_69
timestamp 1669390400
transform 1 0 9072 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1669390400
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1669390400
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1669390400
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1669390400
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_208
timestamp 1669390400
transform 1 0 24640 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1669390400
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1669390400
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1669390400
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1669390400
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1669390400
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1669390400
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1669390400
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_357
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_389
timestamp 1669390400
transform 1 0 44912 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_397
timestamp 1669390400
transform 1 0 45808 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_404
timestamp 1669390400
transform 1 0 46592 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_408
timestamp 1669390400
transform 1 0 47040 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_424
timestamp 1669390400
transform 1 0 48832 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_428
timestamp 1669390400
transform 1 0 49280 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_460
timestamp 1669390400
transform 1 0 52864 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_476
timestamp 1669390400
transform 1 0 54656 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_482
timestamp 1669390400
transform 1 0 55328 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_486
timestamp 1669390400
transform 1 0 55776 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_490
timestamp 1669390400
transform 1 0 56224 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_494
timestamp 1669390400
transform 1 0 56672 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1669390400
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_499
timestamp 1669390400
transform 1 0 57232 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_531
timestamp 1669390400
transform 1 0 60816 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_547
timestamp 1669390400
transform 1 0 62608 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_549
timestamp 1669390400
transform 1 0 62832 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_552
timestamp 1669390400
transform 1 0 63168 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_556
timestamp 1669390400
transform 1 0 63616 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_560
timestamp 1669390400
transform 1 0 64064 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_570
timestamp 1669390400
transform 1 0 65184 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_634
timestamp 1669390400
transform 1 0 72352 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1669390400
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_641
timestamp 1669390400
transform 1 0 73136 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_705
timestamp 1669390400
transform 1 0 80304 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_709
timestamp 1669390400
transform 1 0 80752 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_712
timestamp 1669390400
transform 1 0 81088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_776
timestamp 1669390400
transform 1 0 88256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_780
timestamp 1669390400
transform 1 0 88704 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_783
timestamp 1669390400
transform 1 0 89040 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_847
timestamp 1669390400
transform 1 0 96208 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_851
timestamp 1669390400
transform 1 0 96656 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_854
timestamp 1669390400
transform 1 0 96992 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_918
timestamp 1669390400
transform 1 0 104160 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_922
timestamp 1669390400
transform 1 0 104608 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_925
timestamp 1669390400
transform 1 0 104944 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_989
timestamp 1669390400
transform 1 0 112112 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_993
timestamp 1669390400
transform 1 0 112560 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_996
timestamp 1669390400
transform 1 0 112896 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1004
timestamp 1669390400
transform 1 0 113792 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_1007
timestamp 1669390400
transform 1 0 114128 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_1023
timestamp 1669390400
transform 1 0 115920 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1040
timestamp 1669390400
transform 1 0 117824 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1044
timestamp 1669390400
transform 1 0 118272 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_17
timestamp 1669390400
transform 1 0 3248 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_33
timestamp 1669390400
transform 1 0 5040 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1669390400
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1669390400
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1669390400
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1669390400
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1669390400
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1669390400
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1669390400
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1669390400
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1669390400
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1669390400
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1669390400
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1669390400
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1669390400
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1669390400
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1669390400
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1669390400
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1669390400
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1669390400
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_463
timestamp 1669390400
transform 1 0 53200 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_479
timestamp 1669390400
transform 1 0 54992 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_489
timestamp 1669390400
transform 1 0 56112 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_521
timestamp 1669390400
transform 1 0 59696 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_529
timestamp 1669390400
transform 1 0 60592 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1669390400
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1669390400
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1669390400
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1669390400
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_605
timestamp 1669390400
transform 1 0 69104 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_669
timestamp 1669390400
transform 1 0 76272 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1669390400
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_676
timestamp 1669390400
transform 1 0 77056 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_740
timestamp 1669390400
transform 1 0 84224 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_744
timestamp 1669390400
transform 1 0 84672 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_747
timestamp 1669390400
transform 1 0 85008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_811
timestamp 1669390400
transform 1 0 92176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_815
timestamp 1669390400
transform 1 0 92624 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_818
timestamp 1669390400
transform 1 0 92960 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_882
timestamp 1669390400
transform 1 0 100128 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_886
timestamp 1669390400
transform 1 0 100576 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_889
timestamp 1669390400
transform 1 0 100912 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_953
timestamp 1669390400
transform 1 0 108080 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_957
timestamp 1669390400
transform 1 0 108528 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_960
timestamp 1669390400
transform 1 0 108864 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_992
timestamp 1669390400
transform 1 0 112448 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1008
timestamp 1669390400
transform 1 0 114240 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_1011
timestamp 1669390400
transform 1 0 114576 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_1027
timestamp 1669390400
transform 1 0 116368 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1031
timestamp 1669390400
transform 1 0 116816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_1034
timestamp 1669390400
transform 1 0 117152 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_1042
timestamp 1669390400
transform 1 0 118048 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1044
timestamp 1669390400
transform 1 0 118272 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_6
timestamp 1669390400
transform 1 0 2016 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_8
timestamp 1669390400
transform 1 0 2240 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_15
timestamp 1669390400
transform 1 0 3024 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_19
timestamp 1669390400
transform 1 0 3472 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_51
timestamp 1669390400
transform 1 0 7056 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_67
timestamp 1669390400
transform 1 0 8848 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1669390400
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1669390400
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1669390400
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1669390400
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1669390400
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1669390400
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1669390400
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1669390400
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1669390400
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1669390400
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1669390400
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1669390400
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1669390400
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1669390400
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1669390400
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1669390400
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1669390400
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1669390400
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1669390400
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1669390400
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_570
timestamp 1669390400
transform 1 0 65184 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_634
timestamp 1669390400
transform 1 0 72352 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1669390400
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_641
timestamp 1669390400
transform 1 0 73136 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_705
timestamp 1669390400
transform 1 0 80304 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_709
timestamp 1669390400
transform 1 0 80752 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_712
timestamp 1669390400
transform 1 0 81088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_776
timestamp 1669390400
transform 1 0 88256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_780
timestamp 1669390400
transform 1 0 88704 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_783
timestamp 1669390400
transform 1 0 89040 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_847
timestamp 1669390400
transform 1 0 96208 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_851
timestamp 1669390400
transform 1 0 96656 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_854
timestamp 1669390400
transform 1 0 96992 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_918
timestamp 1669390400
transform 1 0 104160 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_922
timestamp 1669390400
transform 1 0 104608 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_925
timestamp 1669390400
transform 1 0 104944 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_989
timestamp 1669390400
transform 1 0 112112 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_993
timestamp 1669390400
transform 1 0 112560 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_996
timestamp 1669390400
transform 1 0 112896 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1012
timestamp 1669390400
transform 1 0 114688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_1016
timestamp 1669390400
transform 1 0 115136 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1018
timestamp 1669390400
transform 1 0 115360 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_1021
timestamp 1669390400
transform 1 0 115696 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_1025
timestamp 1669390400
transform 1 0 116144 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1041
timestamp 1669390400
transform 1 0 117936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_5
timestamp 1669390400
transform 1 0 1904 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_21
timestamp 1669390400
transform 1 0 3696 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_29
timestamp 1669390400
transform 1 0 4592 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_33
timestamp 1669390400
transform 1 0 5040 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1669390400
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1669390400
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1669390400
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1669390400
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1669390400
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1669390400
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1669390400
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1669390400
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1669390400
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1669390400
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1669390400
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1669390400
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1669390400
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1669390400
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1669390400
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1669390400
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1669390400
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1669390400
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1669390400
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1669390400
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1669390400
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1669390400
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1669390400
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_605
timestamp 1669390400
transform 1 0 69104 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_669
timestamp 1669390400
transform 1 0 76272 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_673
timestamp 1669390400
transform 1 0 76720 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_676
timestamp 1669390400
transform 1 0 77056 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_740
timestamp 1669390400
transform 1 0 84224 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_744
timestamp 1669390400
transform 1 0 84672 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_747
timestamp 1669390400
transform 1 0 85008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_811
timestamp 1669390400
transform 1 0 92176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_815
timestamp 1669390400
transform 1 0 92624 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_818
timestamp 1669390400
transform 1 0 92960 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_882
timestamp 1669390400
transform 1 0 100128 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_886
timestamp 1669390400
transform 1 0 100576 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_889
timestamp 1669390400
transform 1 0 100912 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_953
timestamp 1669390400
transform 1 0 108080 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_957
timestamp 1669390400
transform 1 0 108528 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_960
timestamp 1669390400
transform 1 0 108864 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1024
timestamp 1669390400
transform 1 0 116032 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1028
timestamp 1669390400
transform 1 0 116480 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_1031
timestamp 1669390400
transform 1 0 116816 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1039
timestamp 1669390400
transform 1 0 117712 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1044
timestamp 1669390400
transform 1 0 118272 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_19
timestamp 1669390400
transform 1 0 3472 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_51
timestamp 1669390400
transform 1 0 7056 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_67
timestamp 1669390400
transform 1 0 8848 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1669390400
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1669390400
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1669390400
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1669390400
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1669390400
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1669390400
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1669390400
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1669390400
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1669390400
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1669390400
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1669390400
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1669390400
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1669390400
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1669390400
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1669390400
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1669390400
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1669390400
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1669390400
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1669390400
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1669390400
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_570
timestamp 1669390400
transform 1 0 65184 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_634
timestamp 1669390400
transform 1 0 72352 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1669390400
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_641
timestamp 1669390400
transform 1 0 73136 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_705
timestamp 1669390400
transform 1 0 80304 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_709
timestamp 1669390400
transform 1 0 80752 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_712
timestamp 1669390400
transform 1 0 81088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_776
timestamp 1669390400
transform 1 0 88256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_780
timestamp 1669390400
transform 1 0 88704 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_783
timestamp 1669390400
transform 1 0 89040 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_847
timestamp 1669390400
transform 1 0 96208 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_851
timestamp 1669390400
transform 1 0 96656 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_854
timestamp 1669390400
transform 1 0 96992 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_918
timestamp 1669390400
transform 1 0 104160 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_922
timestamp 1669390400
transform 1 0 104608 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_925
timestamp 1669390400
transform 1 0 104944 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_989
timestamp 1669390400
transform 1 0 112112 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_993
timestamp 1669390400
transform 1 0 112560 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_996
timestamp 1669390400
transform 1 0 112896 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_1028
timestamp 1669390400
transform 1 0 116480 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1044
timestamp 1669390400
transform 1 0 118272 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1669390400
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1669390400
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1669390400
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1669390400
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1669390400
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1669390400
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1669390400
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1669390400
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1669390400
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1669390400
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1669390400
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1669390400
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1669390400
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1669390400
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1669390400
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1669390400
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1669390400
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1669390400
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1669390400
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1669390400
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1669390400
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1669390400
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1669390400
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_598
timestamp 1669390400
transform 1 0 68320 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1669390400
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_605
timestamp 1669390400
transform 1 0 69104 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_669
timestamp 1669390400
transform 1 0 76272 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1669390400
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_676
timestamp 1669390400
transform 1 0 77056 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_740
timestamp 1669390400
transform 1 0 84224 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_744
timestamp 1669390400
transform 1 0 84672 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_747
timestamp 1669390400
transform 1 0 85008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_811
timestamp 1669390400
transform 1 0 92176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_815
timestamp 1669390400
transform 1 0 92624 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_818
timestamp 1669390400
transform 1 0 92960 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_882
timestamp 1669390400
transform 1 0 100128 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_886
timestamp 1669390400
transform 1 0 100576 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_889
timestamp 1669390400
transform 1 0 100912 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_953
timestamp 1669390400
transform 1 0 108080 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_957
timestamp 1669390400
transform 1 0 108528 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_960
timestamp 1669390400
transform 1 0 108864 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1024
timestamp 1669390400
transform 1 0 116032 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1028
timestamp 1669390400
transform 1 0 116480 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_1031
timestamp 1669390400
transform 1 0 116816 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1039
timestamp 1669390400
transform 1 0 117712 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_1043
timestamp 1669390400
transform 1 0 118160 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_66
timestamp 1669390400
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_70
timestamp 1669390400
transform 1 0 9184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1669390400
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1669390400
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1669390400
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1669390400
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1669390400
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1669390400
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1669390400
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1669390400
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1669390400
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1669390400
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1669390400
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1669390400
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1669390400
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1669390400
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1669390400
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1669390400
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1669390400
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1669390400
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1669390400
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_570
timestamp 1669390400
transform 1 0 65184 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_634
timestamp 1669390400
transform 1 0 72352 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1669390400
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_641
timestamp 1669390400
transform 1 0 73136 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_705
timestamp 1669390400
transform 1 0 80304 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_709
timestamp 1669390400
transform 1 0 80752 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_712
timestamp 1669390400
transform 1 0 81088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_776
timestamp 1669390400
transform 1 0 88256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_780
timestamp 1669390400
transform 1 0 88704 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_783
timestamp 1669390400
transform 1 0 89040 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_847
timestamp 1669390400
transform 1 0 96208 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_851
timestamp 1669390400
transform 1 0 96656 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_854
timestamp 1669390400
transform 1 0 96992 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_918
timestamp 1669390400
transform 1 0 104160 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_922
timestamp 1669390400
transform 1 0 104608 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_925
timestamp 1669390400
transform 1 0 104944 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_989
timestamp 1669390400
transform 1 0 112112 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_993
timestamp 1669390400
transform 1 0 112560 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_996
timestamp 1669390400
transform 1 0 112896 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_1028
timestamp 1669390400
transform 1 0 116480 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1044
timestamp 1669390400
transform 1 0 118272 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1669390400
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1669390400
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1669390400
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1669390400
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1669390400
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1669390400
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1669390400
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1669390400
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1669390400
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1669390400
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1669390400
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1669390400
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1669390400
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1669390400
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1669390400
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1669390400
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1669390400
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1669390400
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1669390400
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1669390400
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1669390400
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1669390400
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1669390400
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_605
timestamp 1669390400
transform 1 0 69104 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_669
timestamp 1669390400
transform 1 0 76272 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1669390400
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_676
timestamp 1669390400
transform 1 0 77056 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_740
timestamp 1669390400
transform 1 0 84224 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_744
timestamp 1669390400
transform 1 0 84672 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_747
timestamp 1669390400
transform 1 0 85008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_811
timestamp 1669390400
transform 1 0 92176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_815
timestamp 1669390400
transform 1 0 92624 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_818
timestamp 1669390400
transform 1 0 92960 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_882
timestamp 1669390400
transform 1 0 100128 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_886
timestamp 1669390400
transform 1 0 100576 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_889
timestamp 1669390400
transform 1 0 100912 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_953
timestamp 1669390400
transform 1 0 108080 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_957
timestamp 1669390400
transform 1 0 108528 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_960
timestamp 1669390400
transform 1 0 108864 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_992
timestamp 1669390400
transform 1 0 112448 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1008
timestamp 1669390400
transform 1 0 114240 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1028
timestamp 1669390400
transform 1 0 116480 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1031
timestamp 1669390400
transform 1 0 116816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_1034
timestamp 1669390400
transform 1 0 117152 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_1042
timestamp 1669390400
transform 1 0 118048 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1044
timestamp 1669390400
transform 1 0 118272 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_6
timestamp 1669390400
transform 1 0 2016 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_8
timestamp 1669390400
transform 1 0 2240 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_15
timestamp 1669390400
transform 1 0 3024 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_19
timestamp 1669390400
transform 1 0 3472 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_51
timestamp 1669390400
transform 1 0 7056 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_67
timestamp 1669390400
transform 1 0 8848 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1669390400
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1669390400
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1669390400
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1669390400
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1669390400
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1669390400
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1669390400
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1669390400
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1669390400
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1669390400
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1669390400
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1669390400
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1669390400
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1669390400
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1669390400
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1669390400
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1669390400
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1669390400
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1669390400
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1669390400
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1669390400
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1669390400
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1669390400
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_641
timestamp 1669390400
transform 1 0 73136 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_705
timestamp 1669390400
transform 1 0 80304 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_709
timestamp 1669390400
transform 1 0 80752 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_712
timestamp 1669390400
transform 1 0 81088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_776
timestamp 1669390400
transform 1 0 88256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_780
timestamp 1669390400
transform 1 0 88704 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_783
timestamp 1669390400
transform 1 0 89040 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_847
timestamp 1669390400
transform 1 0 96208 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_851
timestamp 1669390400
transform 1 0 96656 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_854
timestamp 1669390400
transform 1 0 96992 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_918
timestamp 1669390400
transform 1 0 104160 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_922
timestamp 1669390400
transform 1 0 104608 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_925
timestamp 1669390400
transform 1 0 104944 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_989
timestamp 1669390400
transform 1 0 112112 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_993
timestamp 1669390400
transform 1 0 112560 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_996
timestamp 1669390400
transform 1 0 112896 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_1028
timestamp 1669390400
transform 1 0 116480 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1044
timestamp 1669390400
transform 1 0 118272 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_17
timestamp 1669390400
transform 1 0 3248 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_33
timestamp 1669390400
transform 1 0 5040 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1669390400
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1669390400
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1669390400
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1669390400
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1669390400
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1669390400
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1669390400
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1669390400
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1669390400
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1669390400
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1669390400
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1669390400
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1669390400
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1669390400
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1669390400
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1669390400
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_463
timestamp 1669390400
transform 1 0 53200 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1669390400
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1669390400
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1669390400
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1669390400
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1669390400
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_605
timestamp 1669390400
transform 1 0 69104 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_669
timestamp 1669390400
transform 1 0 76272 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_673
timestamp 1669390400
transform 1 0 76720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_676
timestamp 1669390400
transform 1 0 77056 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_740
timestamp 1669390400
transform 1 0 84224 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_744
timestamp 1669390400
transform 1 0 84672 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_747
timestamp 1669390400
transform 1 0 85008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_811
timestamp 1669390400
transform 1 0 92176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_815
timestamp 1669390400
transform 1 0 92624 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_818
timestamp 1669390400
transform 1 0 92960 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_882
timestamp 1669390400
transform 1 0 100128 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_886
timestamp 1669390400
transform 1 0 100576 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_889
timestamp 1669390400
transform 1 0 100912 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_953
timestamp 1669390400
transform 1 0 108080 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_957
timestamp 1669390400
transform 1 0 108528 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_960
timestamp 1669390400
transform 1 0 108864 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_992
timestamp 1669390400
transform 1 0 112448 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1008
timestamp 1669390400
transform 1 0 114240 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_1011
timestamp 1669390400
transform 1 0 114576 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_1027
timestamp 1669390400
transform 1 0 116368 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_1031
timestamp 1669390400
transform 1 0 116816 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1039
timestamp 1669390400
transform 1 0 117712 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_1043
timestamp 1669390400
transform 1 0 118160 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_28
timestamp 1669390400
transform 1 0 4480 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_60
timestamp 1669390400
transform 1 0 8064 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_68
timestamp 1669390400
transform 1 0 8960 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_70
timestamp 1669390400
transform 1 0 9184 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_73
timestamp 1669390400
transform 1 0 9520 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_137
timestamp 1669390400
transform 1 0 16688 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_141
timestamp 1669390400
transform 1 0 17136 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_144
timestamp 1669390400
transform 1 0 17472 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_208
timestamp 1669390400
transform 1 0 24640 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_212
timestamp 1669390400
transform 1 0 25088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_215
timestamp 1669390400
transform 1 0 25424 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_279
timestamp 1669390400
transform 1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_283
timestamp 1669390400
transform 1 0 33040 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_286
timestamp 1669390400
transform 1 0 33376 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_350
timestamp 1669390400
transform 1 0 40544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_354
timestamp 1669390400
transform 1 0 40992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_357
timestamp 1669390400
transform 1 0 41328 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_421
timestamp 1669390400
transform 1 0 48496 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_425
timestamp 1669390400
transform 1 0 48944 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_428
timestamp 1669390400
transform 1 0 49280 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_492
timestamp 1669390400
transform 1 0 56448 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_496
timestamp 1669390400
transform 1 0 56896 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_499
timestamp 1669390400
transform 1 0 57232 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_563
timestamp 1669390400
transform 1 0 64400 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_567
timestamp 1669390400
transform 1 0 64848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_570
timestamp 1669390400
transform 1 0 65184 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_634
timestamp 1669390400
transform 1 0 72352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_638
timestamp 1669390400
transform 1 0 72800 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_641
timestamp 1669390400
transform 1 0 73136 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_705
timestamp 1669390400
transform 1 0 80304 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_709
timestamp 1669390400
transform 1 0 80752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_712
timestamp 1669390400
transform 1 0 81088 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_776
timestamp 1669390400
transform 1 0 88256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_780
timestamp 1669390400
transform 1 0 88704 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_783
timestamp 1669390400
transform 1 0 89040 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_847
timestamp 1669390400
transform 1 0 96208 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_851
timestamp 1669390400
transform 1 0 96656 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_854
timestamp 1669390400
transform 1 0 96992 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_918
timestamp 1669390400
transform 1 0 104160 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_922
timestamp 1669390400
transform 1 0 104608 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_925
timestamp 1669390400
transform 1 0 104944 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_989
timestamp 1669390400
transform 1 0 112112 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_993
timestamp 1669390400
transform 1 0 112560 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_996
timestamp 1669390400
transform 1 0 112896 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_1028
timestamp 1669390400
transform 1 0 116480 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1044
timestamp 1669390400
transform 1 0 118272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_2
timestamp 1669390400
transform 1 0 1568 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_5
timestamp 1669390400
transform 1 0 1904 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_21
timestamp 1669390400
transform 1 0 3696 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_29
timestamp 1669390400
transform 1 0 4592 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_33
timestamp 1669390400
transform 1 0 5040 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_37
timestamp 1669390400
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_101
timestamp 1669390400
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_105
timestamp 1669390400
transform 1 0 13104 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_108
timestamp 1669390400
transform 1 0 13440 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_172
timestamp 1669390400
transform 1 0 20608 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_176
timestamp 1669390400
transform 1 0 21056 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_179
timestamp 1669390400
transform 1 0 21392 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_243
timestamp 1669390400
transform 1 0 28560 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_247
timestamp 1669390400
transform 1 0 29008 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_250
timestamp 1669390400
transform 1 0 29344 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_314
timestamp 1669390400
transform 1 0 36512 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_318
timestamp 1669390400
transform 1 0 36960 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_321
timestamp 1669390400
transform 1 0 37296 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_385
timestamp 1669390400
transform 1 0 44464 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_389
timestamp 1669390400
transform 1 0 44912 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_392
timestamp 1669390400
transform 1 0 45248 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_456
timestamp 1669390400
transform 1 0 52416 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_460
timestamp 1669390400
transform 1 0 52864 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_463
timestamp 1669390400
transform 1 0 53200 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_527
timestamp 1669390400
transform 1 0 60368 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_531
timestamp 1669390400
transform 1 0 60816 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_534
timestamp 1669390400
transform 1 0 61152 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_598
timestamp 1669390400
transform 1 0 68320 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_602
timestamp 1669390400
transform 1 0 68768 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_605
timestamp 1669390400
transform 1 0 69104 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_669
timestamp 1669390400
transform 1 0 76272 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_673
timestamp 1669390400
transform 1 0 76720 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_676
timestamp 1669390400
transform 1 0 77056 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_740
timestamp 1669390400
transform 1 0 84224 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_744
timestamp 1669390400
transform 1 0 84672 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_747
timestamp 1669390400
transform 1 0 85008 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_811
timestamp 1669390400
transform 1 0 92176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_815
timestamp 1669390400
transform 1 0 92624 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_818
timestamp 1669390400
transform 1 0 92960 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_882
timestamp 1669390400
transform 1 0 100128 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_886
timestamp 1669390400
transform 1 0 100576 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_889
timestamp 1669390400
transform 1 0 100912 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_953
timestamp 1669390400
transform 1 0 108080 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_957
timestamp 1669390400
transform 1 0 108528 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_960
timestamp 1669390400
transform 1 0 108864 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1024
timestamp 1669390400
transform 1 0 116032 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1028
timestamp 1669390400
transform 1 0 116480 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_1031
timestamp 1669390400
transform 1 0 116816 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1039
timestamp 1669390400
transform 1 0 117712 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_1043
timestamp 1669390400
transform 1 0 118160 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_2
timestamp 1669390400
transform 1 0 1568 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_66
timestamp 1669390400
transform 1 0 8736 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_70
timestamp 1669390400
transform 1 0 9184 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_73
timestamp 1669390400
transform 1 0 9520 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_137
timestamp 1669390400
transform 1 0 16688 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_141
timestamp 1669390400
transform 1 0 17136 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_144
timestamp 1669390400
transform 1 0 17472 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_208
timestamp 1669390400
transform 1 0 24640 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_212
timestamp 1669390400
transform 1 0 25088 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_215
timestamp 1669390400
transform 1 0 25424 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_279
timestamp 1669390400
transform 1 0 32592 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_283
timestamp 1669390400
transform 1 0 33040 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_286
timestamp 1669390400
transform 1 0 33376 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_350
timestamp 1669390400
transform 1 0 40544 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_354
timestamp 1669390400
transform 1 0 40992 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_357
timestamp 1669390400
transform 1 0 41328 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_421
timestamp 1669390400
transform 1 0 48496 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_425
timestamp 1669390400
transform 1 0 48944 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_428
timestamp 1669390400
transform 1 0 49280 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_492
timestamp 1669390400
transform 1 0 56448 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_496
timestamp 1669390400
transform 1 0 56896 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_499
timestamp 1669390400
transform 1 0 57232 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_563
timestamp 1669390400
transform 1 0 64400 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_567
timestamp 1669390400
transform 1 0 64848 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_570
timestamp 1669390400
transform 1 0 65184 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_634
timestamp 1669390400
transform 1 0 72352 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_638
timestamp 1669390400
transform 1 0 72800 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_641
timestamp 1669390400
transform 1 0 73136 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_705
timestamp 1669390400
transform 1 0 80304 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_709
timestamp 1669390400
transform 1 0 80752 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_712
timestamp 1669390400
transform 1 0 81088 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_776
timestamp 1669390400
transform 1 0 88256 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_780
timestamp 1669390400
transform 1 0 88704 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_783
timestamp 1669390400
transform 1 0 89040 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_847
timestamp 1669390400
transform 1 0 96208 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_851
timestamp 1669390400
transform 1 0 96656 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_854
timestamp 1669390400
transform 1 0 96992 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_918
timestamp 1669390400
transform 1 0 104160 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_922
timestamp 1669390400
transform 1 0 104608 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_925
timestamp 1669390400
transform 1 0 104944 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_989
timestamp 1669390400
transform 1 0 112112 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_993
timestamp 1669390400
transform 1 0 112560 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_996
timestamp 1669390400
transform 1 0 112896 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1012
timestamp 1669390400
transform 1 0 114688 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_1038
timestamp 1669390400
transform 1 0 117600 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_1042
timestamp 1669390400
transform 1 0 118048 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1044
timestamp 1669390400
transform 1 0 118272 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_2
timestamp 1669390400
transform 1 0 1568 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_17
timestamp 1669390400
transform 1 0 3248 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_96_21
timestamp 1669390400
transform 1 0 3696 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_29
timestamp 1669390400
transform 1 0 4592 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_33
timestamp 1669390400
transform 1 0 5040 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_37
timestamp 1669390400
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_101
timestamp 1669390400
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_105
timestamp 1669390400
transform 1 0 13104 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_108
timestamp 1669390400
transform 1 0 13440 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_172
timestamp 1669390400
transform 1 0 20608 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_176
timestamp 1669390400
transform 1 0 21056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_179
timestamp 1669390400
transform 1 0 21392 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_243
timestamp 1669390400
transform 1 0 28560 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_247
timestamp 1669390400
transform 1 0 29008 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_250
timestamp 1669390400
transform 1 0 29344 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_314
timestamp 1669390400
transform 1 0 36512 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_318
timestamp 1669390400
transform 1 0 36960 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_321
timestamp 1669390400
transform 1 0 37296 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_385
timestamp 1669390400
transform 1 0 44464 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_389
timestamp 1669390400
transform 1 0 44912 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_392
timestamp 1669390400
transform 1 0 45248 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_456
timestamp 1669390400
transform 1 0 52416 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_460
timestamp 1669390400
transform 1 0 52864 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_463
timestamp 1669390400
transform 1 0 53200 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_527
timestamp 1669390400
transform 1 0 60368 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_531
timestamp 1669390400
transform 1 0 60816 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_534
timestamp 1669390400
transform 1 0 61152 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_598
timestamp 1669390400
transform 1 0 68320 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_602
timestamp 1669390400
transform 1 0 68768 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_605
timestamp 1669390400
transform 1 0 69104 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_669
timestamp 1669390400
transform 1 0 76272 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_673
timestamp 1669390400
transform 1 0 76720 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_676
timestamp 1669390400
transform 1 0 77056 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_740
timestamp 1669390400
transform 1 0 84224 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_744
timestamp 1669390400
transform 1 0 84672 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_747
timestamp 1669390400
transform 1 0 85008 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_811
timestamp 1669390400
transform 1 0 92176 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_815
timestamp 1669390400
transform 1 0 92624 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_818
timestamp 1669390400
transform 1 0 92960 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_882
timestamp 1669390400
transform 1 0 100128 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_886
timestamp 1669390400
transform 1 0 100576 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_889
timestamp 1669390400
transform 1 0 100912 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_953
timestamp 1669390400
transform 1 0 108080 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_957
timestamp 1669390400
transform 1 0 108528 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_960
timestamp 1669390400
transform 1 0 108864 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1024
timestamp 1669390400
transform 1 0 116032 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1028
timestamp 1669390400
transform 1 0 116480 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_96_1031
timestamp 1669390400
transform 1 0 116816 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1039
timestamp 1669390400
transform 1 0 117712 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1044
timestamp 1669390400
transform 1 0 118272 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_2
timestamp 1669390400
transform 1 0 1568 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_6
timestamp 1669390400
transform 1 0 2016 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_8
timestamp 1669390400
transform 1 0 2240 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_15
timestamp 1669390400
transform 1 0 3024 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_97_19
timestamp 1669390400
transform 1 0 3472 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_51
timestamp 1669390400
transform 1 0 7056 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_67
timestamp 1669390400
transform 1 0 8848 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_73
timestamp 1669390400
transform 1 0 9520 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_137
timestamp 1669390400
transform 1 0 16688 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_141
timestamp 1669390400
transform 1 0 17136 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_144
timestamp 1669390400
transform 1 0 17472 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_208
timestamp 1669390400
transform 1 0 24640 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_212
timestamp 1669390400
transform 1 0 25088 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_215
timestamp 1669390400
transform 1 0 25424 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_279
timestamp 1669390400
transform 1 0 32592 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_283
timestamp 1669390400
transform 1 0 33040 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_286
timestamp 1669390400
transform 1 0 33376 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_350
timestamp 1669390400
transform 1 0 40544 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_354
timestamp 1669390400
transform 1 0 40992 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_357
timestamp 1669390400
transform 1 0 41328 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_421
timestamp 1669390400
transform 1 0 48496 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_425
timestamp 1669390400
transform 1 0 48944 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_428
timestamp 1669390400
transform 1 0 49280 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_492
timestamp 1669390400
transform 1 0 56448 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_496
timestamp 1669390400
transform 1 0 56896 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_499
timestamp 1669390400
transform 1 0 57232 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_563
timestamp 1669390400
transform 1 0 64400 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_567
timestamp 1669390400
transform 1 0 64848 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_570
timestamp 1669390400
transform 1 0 65184 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_634
timestamp 1669390400
transform 1 0 72352 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_638
timestamp 1669390400
transform 1 0 72800 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_641
timestamp 1669390400
transform 1 0 73136 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_705
timestamp 1669390400
transform 1 0 80304 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_709
timestamp 1669390400
transform 1 0 80752 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_712
timestamp 1669390400
transform 1 0 81088 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_776
timestamp 1669390400
transform 1 0 88256 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_780
timestamp 1669390400
transform 1 0 88704 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_783
timestamp 1669390400
transform 1 0 89040 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_847
timestamp 1669390400
transform 1 0 96208 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_851
timestamp 1669390400
transform 1 0 96656 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_854
timestamp 1669390400
transform 1 0 96992 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_918
timestamp 1669390400
transform 1 0 104160 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_922
timestamp 1669390400
transform 1 0 104608 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_925
timestamp 1669390400
transform 1 0 104944 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_989
timestamp 1669390400
transform 1 0 112112 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_993
timestamp 1669390400
transform 1 0 112560 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_996
timestamp 1669390400
transform 1 0 112896 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1012
timestamp 1669390400
transform 1 0 114688 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_1038
timestamp 1669390400
transform 1 0 117600 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_1042
timestamp 1669390400
transform 1 0 118048 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1044
timestamp 1669390400
transform 1 0 118272 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_2
timestamp 1669390400
transform 1 0 1568 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_98_17
timestamp 1669390400
transform 1 0 3248 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_33
timestamp 1669390400
transform 1 0 5040 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_37
timestamp 1669390400
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_101
timestamp 1669390400
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_105
timestamp 1669390400
transform 1 0 13104 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_108
timestamp 1669390400
transform 1 0 13440 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_172
timestamp 1669390400
transform 1 0 20608 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_176
timestamp 1669390400
transform 1 0 21056 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_179
timestamp 1669390400
transform 1 0 21392 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_243
timestamp 1669390400
transform 1 0 28560 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_247
timestamp 1669390400
transform 1 0 29008 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_250
timestamp 1669390400
transform 1 0 29344 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_314
timestamp 1669390400
transform 1 0 36512 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_318
timestamp 1669390400
transform 1 0 36960 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_321
timestamp 1669390400
transform 1 0 37296 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_385
timestamp 1669390400
transform 1 0 44464 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_389
timestamp 1669390400
transform 1 0 44912 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_392
timestamp 1669390400
transform 1 0 45248 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_456
timestamp 1669390400
transform 1 0 52416 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_460
timestamp 1669390400
transform 1 0 52864 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_463
timestamp 1669390400
transform 1 0 53200 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_527
timestamp 1669390400
transform 1 0 60368 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_531
timestamp 1669390400
transform 1 0 60816 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_534
timestamp 1669390400
transform 1 0 61152 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_598
timestamp 1669390400
transform 1 0 68320 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_602
timestamp 1669390400
transform 1 0 68768 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_605
timestamp 1669390400
transform 1 0 69104 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_669
timestamp 1669390400
transform 1 0 76272 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_673
timestamp 1669390400
transform 1 0 76720 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_676
timestamp 1669390400
transform 1 0 77056 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_740
timestamp 1669390400
transform 1 0 84224 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_744
timestamp 1669390400
transform 1 0 84672 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_747
timestamp 1669390400
transform 1 0 85008 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_811
timestamp 1669390400
transform 1 0 92176 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_815
timestamp 1669390400
transform 1 0 92624 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_818
timestamp 1669390400
transform 1 0 92960 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_882
timestamp 1669390400
transform 1 0 100128 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_886
timestamp 1669390400
transform 1 0 100576 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_889
timestamp 1669390400
transform 1 0 100912 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_953
timestamp 1669390400
transform 1 0 108080 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_957
timestamp 1669390400
transform 1 0 108528 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_960
timestamp 1669390400
transform 1 0 108864 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1024
timestamp 1669390400
transform 1 0 116032 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1028
timestamp 1669390400
transform 1 0 116480 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_98_1031
timestamp 1669390400
transform 1 0 116816 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1039
timestamp 1669390400
transform 1 0 117712 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_1043
timestamp 1669390400
transform 1 0 118160 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_2
timestamp 1669390400
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_66
timestamp 1669390400
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_70
timestamp 1669390400
transform 1 0 9184 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_73
timestamp 1669390400
transform 1 0 9520 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_137
timestamp 1669390400
transform 1 0 16688 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_141
timestamp 1669390400
transform 1 0 17136 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_144
timestamp 1669390400
transform 1 0 17472 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_208
timestamp 1669390400
transform 1 0 24640 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_212
timestamp 1669390400
transform 1 0 25088 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_215
timestamp 1669390400
transform 1 0 25424 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_279
timestamp 1669390400
transform 1 0 32592 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_283
timestamp 1669390400
transform 1 0 33040 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_286
timestamp 1669390400
transform 1 0 33376 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_350
timestamp 1669390400
transform 1 0 40544 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_354
timestamp 1669390400
transform 1 0 40992 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_357
timestamp 1669390400
transform 1 0 41328 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_421
timestamp 1669390400
transform 1 0 48496 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_425
timestamp 1669390400
transform 1 0 48944 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_428
timestamp 1669390400
transform 1 0 49280 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_492
timestamp 1669390400
transform 1 0 56448 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_496
timestamp 1669390400
transform 1 0 56896 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_499
timestamp 1669390400
transform 1 0 57232 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_563
timestamp 1669390400
transform 1 0 64400 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_567
timestamp 1669390400
transform 1 0 64848 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_570
timestamp 1669390400
transform 1 0 65184 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_634
timestamp 1669390400
transform 1 0 72352 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_638
timestamp 1669390400
transform 1 0 72800 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_641
timestamp 1669390400
transform 1 0 73136 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_705
timestamp 1669390400
transform 1 0 80304 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_709
timestamp 1669390400
transform 1 0 80752 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_712
timestamp 1669390400
transform 1 0 81088 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_776
timestamp 1669390400
transform 1 0 88256 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_780
timestamp 1669390400
transform 1 0 88704 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_783
timestamp 1669390400
transform 1 0 89040 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_847
timestamp 1669390400
transform 1 0 96208 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_851
timestamp 1669390400
transform 1 0 96656 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_854
timestamp 1669390400
transform 1 0 96992 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_918
timestamp 1669390400
transform 1 0 104160 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_922
timestamp 1669390400
transform 1 0 104608 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_925
timestamp 1669390400
transform 1 0 104944 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_989
timestamp 1669390400
transform 1 0 112112 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_993
timestamp 1669390400
transform 1 0 112560 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_99_996
timestamp 1669390400
transform 1 0 112896 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_1028
timestamp 1669390400
transform 1 0 116480 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1044
timestamp 1669390400
transform 1 0 118272 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_2
timestamp 1669390400
transform 1 0 1568 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_6
timestamp 1669390400
transform 1 0 2016 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_8
timestamp 1669390400
transform 1 0 2240 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_15
timestamp 1669390400
transform 1 0 3024 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_100_19
timestamp 1669390400
transform 1 0 3472 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_37
timestamp 1669390400
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_101
timestamp 1669390400
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_105
timestamp 1669390400
transform 1 0 13104 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_108
timestamp 1669390400
transform 1 0 13440 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_172
timestamp 1669390400
transform 1 0 20608 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_176
timestamp 1669390400
transform 1 0 21056 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_179
timestamp 1669390400
transform 1 0 21392 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_243
timestamp 1669390400
transform 1 0 28560 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_247
timestamp 1669390400
transform 1 0 29008 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_250
timestamp 1669390400
transform 1 0 29344 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_314
timestamp 1669390400
transform 1 0 36512 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_318
timestamp 1669390400
transform 1 0 36960 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_321
timestamp 1669390400
transform 1 0 37296 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_385
timestamp 1669390400
transform 1 0 44464 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_389
timestamp 1669390400
transform 1 0 44912 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_392
timestamp 1669390400
transform 1 0 45248 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_456
timestamp 1669390400
transform 1 0 52416 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_460
timestamp 1669390400
transform 1 0 52864 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_463
timestamp 1669390400
transform 1 0 53200 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_527
timestamp 1669390400
transform 1 0 60368 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_531
timestamp 1669390400
transform 1 0 60816 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_534
timestamp 1669390400
transform 1 0 61152 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_598
timestamp 1669390400
transform 1 0 68320 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_602
timestamp 1669390400
transform 1 0 68768 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_605
timestamp 1669390400
transform 1 0 69104 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_669
timestamp 1669390400
transform 1 0 76272 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_673
timestamp 1669390400
transform 1 0 76720 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_676
timestamp 1669390400
transform 1 0 77056 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_740
timestamp 1669390400
transform 1 0 84224 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_744
timestamp 1669390400
transform 1 0 84672 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_747
timestamp 1669390400
transform 1 0 85008 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_811
timestamp 1669390400
transform 1 0 92176 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_815
timestamp 1669390400
transform 1 0 92624 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_818
timestamp 1669390400
transform 1 0 92960 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_882
timestamp 1669390400
transform 1 0 100128 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_886
timestamp 1669390400
transform 1 0 100576 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_889
timestamp 1669390400
transform 1 0 100912 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_953
timestamp 1669390400
transform 1 0 108080 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_957
timestamp 1669390400
transform 1 0 108528 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_960
timestamp 1669390400
transform 1 0 108864 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1024
timestamp 1669390400
transform 1 0 116032 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1028
timestamp 1669390400
transform 1 0 116480 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_1031
timestamp 1669390400
transform 1 0 116816 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1039
timestamp 1669390400
transform 1 0 117712 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_1043
timestamp 1669390400
transform 1 0 118160 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_2
timestamp 1669390400
transform 1 0 1568 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_101_17
timestamp 1669390400
transform 1 0 3248 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_101_49
timestamp 1669390400
transform 1 0 6832 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_65
timestamp 1669390400
transform 1 0 8624 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_69
timestamp 1669390400
transform 1 0 9072 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_73
timestamp 1669390400
transform 1 0 9520 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_137
timestamp 1669390400
transform 1 0 16688 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_141
timestamp 1669390400
transform 1 0 17136 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_144
timestamp 1669390400
transform 1 0 17472 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_208
timestamp 1669390400
transform 1 0 24640 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_212
timestamp 1669390400
transform 1 0 25088 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_215
timestamp 1669390400
transform 1 0 25424 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_279
timestamp 1669390400
transform 1 0 32592 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_283
timestamp 1669390400
transform 1 0 33040 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_286
timestamp 1669390400
transform 1 0 33376 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_350
timestamp 1669390400
transform 1 0 40544 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_354
timestamp 1669390400
transform 1 0 40992 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_357
timestamp 1669390400
transform 1 0 41328 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_421
timestamp 1669390400
transform 1 0 48496 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_425
timestamp 1669390400
transform 1 0 48944 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_428
timestamp 1669390400
transform 1 0 49280 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_492
timestamp 1669390400
transform 1 0 56448 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_496
timestamp 1669390400
transform 1 0 56896 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_499
timestamp 1669390400
transform 1 0 57232 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_563
timestamp 1669390400
transform 1 0 64400 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_567
timestamp 1669390400
transform 1 0 64848 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_570
timestamp 1669390400
transform 1 0 65184 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_634
timestamp 1669390400
transform 1 0 72352 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_638
timestamp 1669390400
transform 1 0 72800 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_641
timestamp 1669390400
transform 1 0 73136 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_705
timestamp 1669390400
transform 1 0 80304 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_709
timestamp 1669390400
transform 1 0 80752 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_712
timestamp 1669390400
transform 1 0 81088 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_776
timestamp 1669390400
transform 1 0 88256 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_780
timestamp 1669390400
transform 1 0 88704 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_783
timestamp 1669390400
transform 1 0 89040 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_847
timestamp 1669390400
transform 1 0 96208 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_851
timestamp 1669390400
transform 1 0 96656 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_854
timestamp 1669390400
transform 1 0 96992 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_918
timestamp 1669390400
transform 1 0 104160 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_922
timestamp 1669390400
transform 1 0 104608 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_925
timestamp 1669390400
transform 1 0 104944 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_989
timestamp 1669390400
transform 1 0 112112 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_993
timestamp 1669390400
transform 1 0 112560 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_101_996
timestamp 1669390400
transform 1 0 112896 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_1028
timestamp 1669390400
transform 1 0 116480 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_1032
timestamp 1669390400
transform 1 0 116928 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1044
timestamp 1669390400
transform 1 0 118272 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_2
timestamp 1669390400
transform 1 0 1568 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_34
timestamp 1669390400
transform 1 0 5152 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_37
timestamp 1669390400
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_101
timestamp 1669390400
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_105
timestamp 1669390400
transform 1 0 13104 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_108
timestamp 1669390400
transform 1 0 13440 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_172
timestamp 1669390400
transform 1 0 20608 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_176
timestamp 1669390400
transform 1 0 21056 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_179
timestamp 1669390400
transform 1 0 21392 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_243
timestamp 1669390400
transform 1 0 28560 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_247
timestamp 1669390400
transform 1 0 29008 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_250
timestamp 1669390400
transform 1 0 29344 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_314
timestamp 1669390400
transform 1 0 36512 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_318
timestamp 1669390400
transform 1 0 36960 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_321
timestamp 1669390400
transform 1 0 37296 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_385
timestamp 1669390400
transform 1 0 44464 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_389
timestamp 1669390400
transform 1 0 44912 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_392
timestamp 1669390400
transform 1 0 45248 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_456
timestamp 1669390400
transform 1 0 52416 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_460
timestamp 1669390400
transform 1 0 52864 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_463
timestamp 1669390400
transform 1 0 53200 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_527
timestamp 1669390400
transform 1 0 60368 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_531
timestamp 1669390400
transform 1 0 60816 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_534
timestamp 1669390400
transform 1 0 61152 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_598
timestamp 1669390400
transform 1 0 68320 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_602
timestamp 1669390400
transform 1 0 68768 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_605
timestamp 1669390400
transform 1 0 69104 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_669
timestamp 1669390400
transform 1 0 76272 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_673
timestamp 1669390400
transform 1 0 76720 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_676
timestamp 1669390400
transform 1 0 77056 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_740
timestamp 1669390400
transform 1 0 84224 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_744
timestamp 1669390400
transform 1 0 84672 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_747
timestamp 1669390400
transform 1 0 85008 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_811
timestamp 1669390400
transform 1 0 92176 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_815
timestamp 1669390400
transform 1 0 92624 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_818
timestamp 1669390400
transform 1 0 92960 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_882
timestamp 1669390400
transform 1 0 100128 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_886
timestamp 1669390400
transform 1 0 100576 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_889
timestamp 1669390400
transform 1 0 100912 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_953
timestamp 1669390400
transform 1 0 108080 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_957
timestamp 1669390400
transform 1 0 108528 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_960
timestamp 1669390400
transform 1 0 108864 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_992
timestamp 1669390400
transform 1 0 112448 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1008
timestamp 1669390400
transform 1 0 114240 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1012
timestamp 1669390400
transform 1 0 114688 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_1027
timestamp 1669390400
transform 1 0 116368 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1031
timestamp 1669390400
transform 1 0 116816 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1038
timestamp 1669390400
transform 1 0 117600 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_1042
timestamp 1669390400
transform 1 0 118048 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1044
timestamp 1669390400
transform 1 0 118272 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_2
timestamp 1669390400
transform 1 0 1568 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_7
timestamp 1669390400
transform 1 0 2128 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_73
timestamp 1669390400
transform 1 0 9520 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_137
timestamp 1669390400
transform 1 0 16688 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_141
timestamp 1669390400
transform 1 0 17136 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_144
timestamp 1669390400
transform 1 0 17472 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_208
timestamp 1669390400
transform 1 0 24640 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_212
timestamp 1669390400
transform 1 0 25088 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_215
timestamp 1669390400
transform 1 0 25424 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_279
timestamp 1669390400
transform 1 0 32592 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_283
timestamp 1669390400
transform 1 0 33040 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_286
timestamp 1669390400
transform 1 0 33376 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_350
timestamp 1669390400
transform 1 0 40544 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_354
timestamp 1669390400
transform 1 0 40992 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_357
timestamp 1669390400
transform 1 0 41328 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_421
timestamp 1669390400
transform 1 0 48496 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_425
timestamp 1669390400
transform 1 0 48944 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_428
timestamp 1669390400
transform 1 0 49280 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_492
timestamp 1669390400
transform 1 0 56448 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_496
timestamp 1669390400
transform 1 0 56896 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_499
timestamp 1669390400
transform 1 0 57232 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_563
timestamp 1669390400
transform 1 0 64400 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_567
timestamp 1669390400
transform 1 0 64848 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_570
timestamp 1669390400
transform 1 0 65184 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_634
timestamp 1669390400
transform 1 0 72352 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_638
timestamp 1669390400
transform 1 0 72800 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_641
timestamp 1669390400
transform 1 0 73136 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_705
timestamp 1669390400
transform 1 0 80304 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_709
timestamp 1669390400
transform 1 0 80752 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_712
timestamp 1669390400
transform 1 0 81088 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_776
timestamp 1669390400
transform 1 0 88256 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_780
timestamp 1669390400
transform 1 0 88704 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_783
timestamp 1669390400
transform 1 0 89040 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_847
timestamp 1669390400
transform 1 0 96208 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_851
timestamp 1669390400
transform 1 0 96656 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_854
timestamp 1669390400
transform 1 0 96992 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_918
timestamp 1669390400
transform 1 0 104160 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_922
timestamp 1669390400
transform 1 0 104608 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_925
timestamp 1669390400
transform 1 0 104944 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_989
timestamp 1669390400
transform 1 0 112112 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_993
timestamp 1669390400
transform 1 0 112560 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_103_996
timestamp 1669390400
transform 1 0 112896 0 -1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_103_1028
timestamp 1669390400
transform 1 0 116480 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1044
timestamp 1669390400
transform 1 0 118272 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_2
timestamp 1669390400
transform 1 0 1568 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_34
timestamp 1669390400
transform 1 0 5152 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_37
timestamp 1669390400
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_101
timestamp 1669390400
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_105
timestamp 1669390400
transform 1 0 13104 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_108
timestamp 1669390400
transform 1 0 13440 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_172
timestamp 1669390400
transform 1 0 20608 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_176
timestamp 1669390400
transform 1 0 21056 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_179
timestamp 1669390400
transform 1 0 21392 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_243
timestamp 1669390400
transform 1 0 28560 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_247
timestamp 1669390400
transform 1 0 29008 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_250
timestamp 1669390400
transform 1 0 29344 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_314
timestamp 1669390400
transform 1 0 36512 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_318
timestamp 1669390400
transform 1 0 36960 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_321
timestamp 1669390400
transform 1 0 37296 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_385
timestamp 1669390400
transform 1 0 44464 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_389
timestamp 1669390400
transform 1 0 44912 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_392
timestamp 1669390400
transform 1 0 45248 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_456
timestamp 1669390400
transform 1 0 52416 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_460
timestamp 1669390400
transform 1 0 52864 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_463
timestamp 1669390400
transform 1 0 53200 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_527
timestamp 1669390400
transform 1 0 60368 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_531
timestamp 1669390400
transform 1 0 60816 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_534
timestamp 1669390400
transform 1 0 61152 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_598
timestamp 1669390400
transform 1 0 68320 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_602
timestamp 1669390400
transform 1 0 68768 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_605
timestamp 1669390400
transform 1 0 69104 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_637
timestamp 1669390400
transform 1 0 72688 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_653
timestamp 1669390400
transform 1 0 74480 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_661
timestamp 1669390400
transform 1 0 75376 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_665
timestamp 1669390400
transform 1 0 75824 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_673
timestamp 1669390400
transform 1 0 76720 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_676
timestamp 1669390400
transform 1 0 77056 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_740
timestamp 1669390400
transform 1 0 84224 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_744
timestamp 1669390400
transform 1 0 84672 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_747
timestamp 1669390400
transform 1 0 85008 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_811
timestamp 1669390400
transform 1 0 92176 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_815
timestamp 1669390400
transform 1 0 92624 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_818
timestamp 1669390400
transform 1 0 92960 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_882
timestamp 1669390400
transform 1 0 100128 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_886
timestamp 1669390400
transform 1 0 100576 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_889
timestamp 1669390400
transform 1 0 100912 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_953
timestamp 1669390400
transform 1 0 108080 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_957
timestamp 1669390400
transform 1 0 108528 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_960
timestamp 1669390400
transform 1 0 108864 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_992
timestamp 1669390400
transform 1 0 112448 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1008
timestamp 1669390400
transform 1 0 114240 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_1011
timestamp 1669390400
transform 1 0 114576 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_1027
timestamp 1669390400
transform 1 0 116368 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_1031
timestamp 1669390400
transform 1 0 116816 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1039
timestamp 1669390400
transform 1 0 117712 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_1043
timestamp 1669390400
transform 1 0 118160 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_2
timestamp 1669390400
transform 1 0 1568 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_7
timestamp 1669390400
transform 1 0 2128 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_73
timestamp 1669390400
transform 1 0 9520 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_137
timestamp 1669390400
transform 1 0 16688 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_141
timestamp 1669390400
transform 1 0 17136 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_144
timestamp 1669390400
transform 1 0 17472 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_208
timestamp 1669390400
transform 1 0 24640 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_212
timestamp 1669390400
transform 1 0 25088 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_215
timestamp 1669390400
transform 1 0 25424 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_279
timestamp 1669390400
transform 1 0 32592 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_283
timestamp 1669390400
transform 1 0 33040 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_286
timestamp 1669390400
transform 1 0 33376 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_350
timestamp 1669390400
transform 1 0 40544 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_354
timestamp 1669390400
transform 1 0 40992 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_357
timestamp 1669390400
transform 1 0 41328 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_421
timestamp 1669390400
transform 1 0 48496 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_425
timestamp 1669390400
transform 1 0 48944 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_428
timestamp 1669390400
transform 1 0 49280 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_492
timestamp 1669390400
transform 1 0 56448 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_496
timestamp 1669390400
transform 1 0 56896 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_499
timestamp 1669390400
transform 1 0 57232 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_563
timestamp 1669390400
transform 1 0 64400 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_567
timestamp 1669390400
transform 1 0 64848 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_570
timestamp 1669390400
transform 1 0 65184 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_634
timestamp 1669390400
transform 1 0 72352 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_638
timestamp 1669390400
transform 1 0 72800 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_641
timestamp 1669390400
transform 1 0 73136 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_705
timestamp 1669390400
transform 1 0 80304 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_709
timestamp 1669390400
transform 1 0 80752 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_712
timestamp 1669390400
transform 1 0 81088 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_776
timestamp 1669390400
transform 1 0 88256 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_780
timestamp 1669390400
transform 1 0 88704 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_783
timestamp 1669390400
transform 1 0 89040 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_847
timestamp 1669390400
transform 1 0 96208 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_851
timestamp 1669390400
transform 1 0 96656 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_854
timestamp 1669390400
transform 1 0 96992 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_918
timestamp 1669390400
transform 1 0 104160 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_922
timestamp 1669390400
transform 1 0 104608 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_925
timestamp 1669390400
transform 1 0 104944 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_989
timestamp 1669390400
transform 1 0 112112 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_993
timestamp 1669390400
transform 1 0 112560 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_105_996
timestamp 1669390400
transform 1 0 112896 0 -1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_105_1028
timestamp 1669390400
transform 1 0 116480 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1044
timestamp 1669390400
transform 1 0 118272 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_2
timestamp 1669390400
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_34
timestamp 1669390400
transform 1 0 5152 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_37
timestamp 1669390400
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_101
timestamp 1669390400
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_105
timestamp 1669390400
transform 1 0 13104 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_108
timestamp 1669390400
transform 1 0 13440 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_172
timestamp 1669390400
transform 1 0 20608 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_176
timestamp 1669390400
transform 1 0 21056 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_179
timestamp 1669390400
transform 1 0 21392 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_243
timestamp 1669390400
transform 1 0 28560 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_247
timestamp 1669390400
transform 1 0 29008 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_250
timestamp 1669390400
transform 1 0 29344 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_314
timestamp 1669390400
transform 1 0 36512 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_318
timestamp 1669390400
transform 1 0 36960 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_321
timestamp 1669390400
transform 1 0 37296 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_385
timestamp 1669390400
transform 1 0 44464 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_389
timestamp 1669390400
transform 1 0 44912 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_392
timestamp 1669390400
transform 1 0 45248 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_456
timestamp 1669390400
transform 1 0 52416 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_460
timestamp 1669390400
transform 1 0 52864 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_463
timestamp 1669390400
transform 1 0 53200 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_527
timestamp 1669390400
transform 1 0 60368 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_531
timestamp 1669390400
transform 1 0 60816 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_534
timestamp 1669390400
transform 1 0 61152 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_598
timestamp 1669390400
transform 1 0 68320 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_602
timestamp 1669390400
transform 1 0 68768 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_605
timestamp 1669390400
transform 1 0 69104 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_669
timestamp 1669390400
transform 1 0 76272 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_673
timestamp 1669390400
transform 1 0 76720 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_676
timestamp 1669390400
transform 1 0 77056 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_740
timestamp 1669390400
transform 1 0 84224 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_744
timestamp 1669390400
transform 1 0 84672 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_747
timestamp 1669390400
transform 1 0 85008 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_811
timestamp 1669390400
transform 1 0 92176 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_815
timestamp 1669390400
transform 1 0 92624 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_818
timestamp 1669390400
transform 1 0 92960 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_882
timestamp 1669390400
transform 1 0 100128 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_886
timestamp 1669390400
transform 1 0 100576 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_889
timestamp 1669390400
transform 1 0 100912 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_953
timestamp 1669390400
transform 1 0 108080 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_957
timestamp 1669390400
transform 1 0 108528 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_960
timestamp 1669390400
transform 1 0 108864 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_992
timestamp 1669390400
transform 1 0 112448 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1008
timestamp 1669390400
transform 1 0 114240 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_1011
timestamp 1669390400
transform 1 0 114576 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_1027
timestamp 1669390400
transform 1 0 116368 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_1031
timestamp 1669390400
transform 1 0 116816 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1039
timestamp 1669390400
transform 1 0 117712 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_1043
timestamp 1669390400
transform 1 0 118160 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_2
timestamp 1669390400
transform 1 0 1568 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_5
timestamp 1669390400
transform 1 0 1904 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_69
timestamp 1669390400
transform 1 0 9072 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_73
timestamp 1669390400
transform 1 0 9520 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_137
timestamp 1669390400
transform 1 0 16688 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_141
timestamp 1669390400
transform 1 0 17136 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_144
timestamp 1669390400
transform 1 0 17472 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_208
timestamp 1669390400
transform 1 0 24640 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_212
timestamp 1669390400
transform 1 0 25088 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_215
timestamp 1669390400
transform 1 0 25424 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_279
timestamp 1669390400
transform 1 0 32592 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_283
timestamp 1669390400
transform 1 0 33040 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_286
timestamp 1669390400
transform 1 0 33376 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_350
timestamp 1669390400
transform 1 0 40544 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_354
timestamp 1669390400
transform 1 0 40992 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_357
timestamp 1669390400
transform 1 0 41328 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_421
timestamp 1669390400
transform 1 0 48496 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_425
timestamp 1669390400
transform 1 0 48944 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_428
timestamp 1669390400
transform 1 0 49280 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_492
timestamp 1669390400
transform 1 0 56448 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_496
timestamp 1669390400
transform 1 0 56896 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_499
timestamp 1669390400
transform 1 0 57232 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_563
timestamp 1669390400
transform 1 0 64400 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_567
timestamp 1669390400
transform 1 0 64848 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_570
timestamp 1669390400
transform 1 0 65184 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_634
timestamp 1669390400
transform 1 0 72352 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_638
timestamp 1669390400
transform 1 0 72800 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_641
timestamp 1669390400
transform 1 0 73136 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_705
timestamp 1669390400
transform 1 0 80304 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_709
timestamp 1669390400
transform 1 0 80752 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_712
timestamp 1669390400
transform 1 0 81088 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_776
timestamp 1669390400
transform 1 0 88256 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_780
timestamp 1669390400
transform 1 0 88704 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_783
timestamp 1669390400
transform 1 0 89040 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_847
timestamp 1669390400
transform 1 0 96208 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_851
timestamp 1669390400
transform 1 0 96656 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_854
timestamp 1669390400
transform 1 0 96992 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_918
timestamp 1669390400
transform 1 0 104160 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_922
timestamp 1669390400
transform 1 0 104608 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_925
timestamp 1669390400
transform 1 0 104944 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_989
timestamp 1669390400
transform 1 0 112112 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_993
timestamp 1669390400
transform 1 0 112560 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_996
timestamp 1669390400
transform 1 0 112896 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1012
timestamp 1669390400
transform 1 0 114688 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_1029
timestamp 1669390400
transform 1 0 116592 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_1033
timestamp 1669390400
transform 1 0 117040 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1041
timestamp 1669390400
transform 1 0 117936 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_2
timestamp 1669390400
transform 1 0 1568 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_19
timestamp 1669390400
transform 1 0 3472 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_37
timestamp 1669390400
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_101
timestamp 1669390400
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_105
timestamp 1669390400
transform 1 0 13104 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_108
timestamp 1669390400
transform 1 0 13440 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_172
timestamp 1669390400
transform 1 0 20608 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_176
timestamp 1669390400
transform 1 0 21056 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_179
timestamp 1669390400
transform 1 0 21392 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_243
timestamp 1669390400
transform 1 0 28560 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_247
timestamp 1669390400
transform 1 0 29008 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_250
timestamp 1669390400
transform 1 0 29344 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_314
timestamp 1669390400
transform 1 0 36512 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_318
timestamp 1669390400
transform 1 0 36960 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_321
timestamp 1669390400
transform 1 0 37296 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_385
timestamp 1669390400
transform 1 0 44464 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_389
timestamp 1669390400
transform 1 0 44912 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_392
timestamp 1669390400
transform 1 0 45248 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_456
timestamp 1669390400
transform 1 0 52416 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_460
timestamp 1669390400
transform 1 0 52864 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_463
timestamp 1669390400
transform 1 0 53200 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_527
timestamp 1669390400
transform 1 0 60368 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_531
timestamp 1669390400
transform 1 0 60816 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_534
timestamp 1669390400
transform 1 0 61152 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_598
timestamp 1669390400
transform 1 0 68320 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_602
timestamp 1669390400
transform 1 0 68768 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_605
timestamp 1669390400
transform 1 0 69104 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_669
timestamp 1669390400
transform 1 0 76272 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_673
timestamp 1669390400
transform 1 0 76720 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_676
timestamp 1669390400
transform 1 0 77056 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_740
timestamp 1669390400
transform 1 0 84224 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_744
timestamp 1669390400
transform 1 0 84672 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_747
timestamp 1669390400
transform 1 0 85008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_811
timestamp 1669390400
transform 1 0 92176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_815
timestamp 1669390400
transform 1 0 92624 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_818
timestamp 1669390400
transform 1 0 92960 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_882
timestamp 1669390400
transform 1 0 100128 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_886
timestamp 1669390400
transform 1 0 100576 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_889
timestamp 1669390400
transform 1 0 100912 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_953
timestamp 1669390400
transform 1 0 108080 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_957
timestamp 1669390400
transform 1 0 108528 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_960
timestamp 1669390400
transform 1 0 108864 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1024
timestamp 1669390400
transform 1 0 116032 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1028
timestamp 1669390400
transform 1 0 116480 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_1031
timestamp 1669390400
transform 1 0 116816 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1039
timestamp 1669390400
transform 1 0 117712 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_1043
timestamp 1669390400
transform 1 0 118160 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_2
timestamp 1669390400
transform 1 0 1568 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_17
timestamp 1669390400
transform 1 0 3248 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_109_21
timestamp 1669390400
transform 1 0 3696 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_53
timestamp 1669390400
transform 1 0 7280 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_69
timestamp 1669390400
transform 1 0 9072 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_73
timestamp 1669390400
transform 1 0 9520 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_137
timestamp 1669390400
transform 1 0 16688 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_141
timestamp 1669390400
transform 1 0 17136 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_144
timestamp 1669390400
transform 1 0 17472 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_208
timestamp 1669390400
transform 1 0 24640 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_212
timestamp 1669390400
transform 1 0 25088 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_215
timestamp 1669390400
transform 1 0 25424 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_279
timestamp 1669390400
transform 1 0 32592 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_283
timestamp 1669390400
transform 1 0 33040 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_286
timestamp 1669390400
transform 1 0 33376 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_350
timestamp 1669390400
transform 1 0 40544 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_354
timestamp 1669390400
transform 1 0 40992 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_357
timestamp 1669390400
transform 1 0 41328 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_421
timestamp 1669390400
transform 1 0 48496 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_425
timestamp 1669390400
transform 1 0 48944 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_428
timestamp 1669390400
transform 1 0 49280 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_492
timestamp 1669390400
transform 1 0 56448 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_496
timestamp 1669390400
transform 1 0 56896 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_499
timestamp 1669390400
transform 1 0 57232 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_563
timestamp 1669390400
transform 1 0 64400 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_567
timestamp 1669390400
transform 1 0 64848 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_570
timestamp 1669390400
transform 1 0 65184 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_634
timestamp 1669390400
transform 1 0 72352 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_638
timestamp 1669390400
transform 1 0 72800 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_641
timestamp 1669390400
transform 1 0 73136 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_705
timestamp 1669390400
transform 1 0 80304 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_709
timestamp 1669390400
transform 1 0 80752 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_712
timestamp 1669390400
transform 1 0 81088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_776
timestamp 1669390400
transform 1 0 88256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_780
timestamp 1669390400
transform 1 0 88704 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_783
timestamp 1669390400
transform 1 0 89040 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_847
timestamp 1669390400
transform 1 0 96208 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_851
timestamp 1669390400
transform 1 0 96656 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_854
timestamp 1669390400
transform 1 0 96992 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_918
timestamp 1669390400
transform 1 0 104160 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_922
timestamp 1669390400
transform 1 0 104608 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_925
timestamp 1669390400
transform 1 0 104944 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_989
timestamp 1669390400
transform 1 0 112112 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_993
timestamp 1669390400
transform 1 0 112560 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_109_996
timestamp 1669390400
transform 1 0 112896 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_1028
timestamp 1669390400
transform 1 0 116480 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1044
timestamp 1669390400
transform 1 0 118272 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_2
timestamp 1669390400
transform 1 0 1568 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_6
timestamp 1669390400
transform 1 0 2016 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_8
timestamp 1669390400
transform 1 0 2240 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_15
timestamp 1669390400
transform 1 0 3024 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_19
timestamp 1669390400
transform 1 0 3472 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_37
timestamp 1669390400
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_101
timestamp 1669390400
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_105
timestamp 1669390400
transform 1 0 13104 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_108
timestamp 1669390400
transform 1 0 13440 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_172
timestamp 1669390400
transform 1 0 20608 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_176
timestamp 1669390400
transform 1 0 21056 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_179
timestamp 1669390400
transform 1 0 21392 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_243
timestamp 1669390400
transform 1 0 28560 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_247
timestamp 1669390400
transform 1 0 29008 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_250
timestamp 1669390400
transform 1 0 29344 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_314
timestamp 1669390400
transform 1 0 36512 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_318
timestamp 1669390400
transform 1 0 36960 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_321
timestamp 1669390400
transform 1 0 37296 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_385
timestamp 1669390400
transform 1 0 44464 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_389
timestamp 1669390400
transform 1 0 44912 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_392
timestamp 1669390400
transform 1 0 45248 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_456
timestamp 1669390400
transform 1 0 52416 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_460
timestamp 1669390400
transform 1 0 52864 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_463
timestamp 1669390400
transform 1 0 53200 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_495
timestamp 1669390400
transform 1 0 56784 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_511
timestamp 1669390400
transform 1 0 58576 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_518
timestamp 1669390400
transform 1 0 59360 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_522
timestamp 1669390400
transform 1 0 59808 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_530
timestamp 1669390400
transform 1 0 60704 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_534
timestamp 1669390400
transform 1 0 61152 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_598
timestamp 1669390400
transform 1 0 68320 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_602
timestamp 1669390400
transform 1 0 68768 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_605
timestamp 1669390400
transform 1 0 69104 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_669
timestamp 1669390400
transform 1 0 76272 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_673
timestamp 1669390400
transform 1 0 76720 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_676
timestamp 1669390400
transform 1 0 77056 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_740
timestamp 1669390400
transform 1 0 84224 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_744
timestamp 1669390400
transform 1 0 84672 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_747
timestamp 1669390400
transform 1 0 85008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_811
timestamp 1669390400
transform 1 0 92176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_815
timestamp 1669390400
transform 1 0 92624 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_818
timestamp 1669390400
transform 1 0 92960 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_882
timestamp 1669390400
transform 1 0 100128 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_886
timestamp 1669390400
transform 1 0 100576 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_889
timestamp 1669390400
transform 1 0 100912 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_953
timestamp 1669390400
transform 1 0 108080 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_957
timestamp 1669390400
transform 1 0 108528 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_960
timestamp 1669390400
transform 1 0 108864 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_992
timestamp 1669390400
transform 1 0 112448 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1008
timestamp 1669390400
transform 1 0 114240 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1012
timestamp 1669390400
transform 1 0 114688 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_1027
timestamp 1669390400
transform 1 0 116368 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1031
timestamp 1669390400
transform 1 0 116816 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_1034
timestamp 1669390400
transform 1 0 117152 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_1042
timestamp 1669390400
transform 1 0 118048 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1044
timestamp 1669390400
transform 1 0 118272 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_2
timestamp 1669390400
transform 1 0 1568 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_111_17
timestamp 1669390400
transform 1 0 3248 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_49
timestamp 1669390400
transform 1 0 6832 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_65
timestamp 1669390400
transform 1 0 8624 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_111_69
timestamp 1669390400
transform 1 0 9072 0 -1 90944
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_73
timestamp 1669390400
transform 1 0 9520 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_137
timestamp 1669390400
transform 1 0 16688 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_141
timestamp 1669390400
transform 1 0 17136 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_144
timestamp 1669390400
transform 1 0 17472 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_208
timestamp 1669390400
transform 1 0 24640 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_212
timestamp 1669390400
transform 1 0 25088 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_215
timestamp 1669390400
transform 1 0 25424 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_279
timestamp 1669390400
transform 1 0 32592 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_283
timestamp 1669390400
transform 1 0 33040 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_286
timestamp 1669390400
transform 1 0 33376 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_350
timestamp 1669390400
transform 1 0 40544 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_354
timestamp 1669390400
transform 1 0 40992 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_357
timestamp 1669390400
transform 1 0 41328 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_421
timestamp 1669390400
transform 1 0 48496 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_425
timestamp 1669390400
transform 1 0 48944 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_428
timestamp 1669390400
transform 1 0 49280 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_492
timestamp 1669390400
transform 1 0 56448 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_496
timestamp 1669390400
transform 1 0 56896 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_499
timestamp 1669390400
transform 1 0 57232 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_563
timestamp 1669390400
transform 1 0 64400 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_567
timestamp 1669390400
transform 1 0 64848 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_570
timestamp 1669390400
transform 1 0 65184 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_634
timestamp 1669390400
transform 1 0 72352 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_638
timestamp 1669390400
transform 1 0 72800 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_641
timestamp 1669390400
transform 1 0 73136 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_705
timestamp 1669390400
transform 1 0 80304 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_709
timestamp 1669390400
transform 1 0 80752 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_712
timestamp 1669390400
transform 1 0 81088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_776
timestamp 1669390400
transform 1 0 88256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_780
timestamp 1669390400
transform 1 0 88704 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_783
timestamp 1669390400
transform 1 0 89040 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_847
timestamp 1669390400
transform 1 0 96208 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_851
timestamp 1669390400
transform 1 0 96656 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_854
timestamp 1669390400
transform 1 0 96992 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_918
timestamp 1669390400
transform 1 0 104160 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_922
timestamp 1669390400
transform 1 0 104608 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_925
timestamp 1669390400
transform 1 0 104944 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_989
timestamp 1669390400
transform 1 0 112112 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_993
timestamp 1669390400
transform 1 0 112560 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_111_996
timestamp 1669390400
transform 1 0 112896 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_1028
timestamp 1669390400
transform 1 0 116480 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1044
timestamp 1669390400
transform 1 0 118272 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_2
timestamp 1669390400
transform 1 0 1568 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_34
timestamp 1669390400
transform 1 0 5152 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_37
timestamp 1669390400
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_101
timestamp 1669390400
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_105
timestamp 1669390400
transform 1 0 13104 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_108
timestamp 1669390400
transform 1 0 13440 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_172
timestamp 1669390400
transform 1 0 20608 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_176
timestamp 1669390400
transform 1 0 21056 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_179
timestamp 1669390400
transform 1 0 21392 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_243
timestamp 1669390400
transform 1 0 28560 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_247
timestamp 1669390400
transform 1 0 29008 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_250
timestamp 1669390400
transform 1 0 29344 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_314
timestamp 1669390400
transform 1 0 36512 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_318
timestamp 1669390400
transform 1 0 36960 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_321
timestamp 1669390400
transform 1 0 37296 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_385
timestamp 1669390400
transform 1 0 44464 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_389
timestamp 1669390400
transform 1 0 44912 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_392
timestamp 1669390400
transform 1 0 45248 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_456
timestamp 1669390400
transform 1 0 52416 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_460
timestamp 1669390400
transform 1 0 52864 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_463
timestamp 1669390400
transform 1 0 53200 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_527
timestamp 1669390400
transform 1 0 60368 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_531
timestamp 1669390400
transform 1 0 60816 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_534
timestamp 1669390400
transform 1 0 61152 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_598
timestamp 1669390400
transform 1 0 68320 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_602
timestamp 1669390400
transform 1 0 68768 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_605
timestamp 1669390400
transform 1 0 69104 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_669
timestamp 1669390400
transform 1 0 76272 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_673
timestamp 1669390400
transform 1 0 76720 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_676
timestamp 1669390400
transform 1 0 77056 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_740
timestamp 1669390400
transform 1 0 84224 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_744
timestamp 1669390400
transform 1 0 84672 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_747
timestamp 1669390400
transform 1 0 85008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_811
timestamp 1669390400
transform 1 0 92176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_815
timestamp 1669390400
transform 1 0 92624 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_818
timestamp 1669390400
transform 1 0 92960 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_882
timestamp 1669390400
transform 1 0 100128 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_886
timestamp 1669390400
transform 1 0 100576 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_889
timestamp 1669390400
transform 1 0 100912 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_953
timestamp 1669390400
transform 1 0 108080 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_957
timestamp 1669390400
transform 1 0 108528 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_960
timestamp 1669390400
transform 1 0 108864 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1024
timestamp 1669390400
transform 1 0 116032 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1028
timestamp 1669390400
transform 1 0 116480 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_1031
timestamp 1669390400
transform 1 0 116816 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1039
timestamp 1669390400
transform 1 0 117712 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_112_1043
timestamp 1669390400
transform 1 0 118160 0 1 90944
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_2
timestamp 1669390400
transform 1 0 1568 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_5
timestamp 1669390400
transform 1 0 1904 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_69
timestamp 1669390400
transform 1 0 9072 0 -1 92512
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_73
timestamp 1669390400
transform 1 0 9520 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_137
timestamp 1669390400
transform 1 0 16688 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_141
timestamp 1669390400
transform 1 0 17136 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_144
timestamp 1669390400
transform 1 0 17472 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_208
timestamp 1669390400
transform 1 0 24640 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_212
timestamp 1669390400
transform 1 0 25088 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_215
timestamp 1669390400
transform 1 0 25424 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_279
timestamp 1669390400
transform 1 0 32592 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_283
timestamp 1669390400
transform 1 0 33040 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_286
timestamp 1669390400
transform 1 0 33376 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_350
timestamp 1669390400
transform 1 0 40544 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_354
timestamp 1669390400
transform 1 0 40992 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_357
timestamp 1669390400
transform 1 0 41328 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_421
timestamp 1669390400
transform 1 0 48496 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_425
timestamp 1669390400
transform 1 0 48944 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_428
timestamp 1669390400
transform 1 0 49280 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_492
timestamp 1669390400
transform 1 0 56448 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_496
timestamp 1669390400
transform 1 0 56896 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_499
timestamp 1669390400
transform 1 0 57232 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_563
timestamp 1669390400
transform 1 0 64400 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_567
timestamp 1669390400
transform 1 0 64848 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_570
timestamp 1669390400
transform 1 0 65184 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_634
timestamp 1669390400
transform 1 0 72352 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_638
timestamp 1669390400
transform 1 0 72800 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_641
timestamp 1669390400
transform 1 0 73136 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_705
timestamp 1669390400
transform 1 0 80304 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_709
timestamp 1669390400
transform 1 0 80752 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_712
timestamp 1669390400
transform 1 0 81088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_776
timestamp 1669390400
transform 1 0 88256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_780
timestamp 1669390400
transform 1 0 88704 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_783
timestamp 1669390400
transform 1 0 89040 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_847
timestamp 1669390400
transform 1 0 96208 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_851
timestamp 1669390400
transform 1 0 96656 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_854
timestamp 1669390400
transform 1 0 96992 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_918
timestamp 1669390400
transform 1 0 104160 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_922
timestamp 1669390400
transform 1 0 104608 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_925
timestamp 1669390400
transform 1 0 104944 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_989
timestamp 1669390400
transform 1 0 112112 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_993
timestamp 1669390400
transform 1 0 112560 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_113_996
timestamp 1669390400
transform 1 0 112896 0 -1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_113_1028
timestamp 1669390400
transform 1 0 116480 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1044
timestamp 1669390400
transform 1 0 118272 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_2
timestamp 1669390400
transform 1 0 1568 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_19
timestamp 1669390400
transform 1 0 3472 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_37
timestamp 1669390400
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_101
timestamp 1669390400
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_105
timestamp 1669390400
transform 1 0 13104 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_108
timestamp 1669390400
transform 1 0 13440 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_172
timestamp 1669390400
transform 1 0 20608 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_176
timestamp 1669390400
transform 1 0 21056 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_179
timestamp 1669390400
transform 1 0 21392 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_243
timestamp 1669390400
transform 1 0 28560 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_247
timestamp 1669390400
transform 1 0 29008 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_250
timestamp 1669390400
transform 1 0 29344 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_314
timestamp 1669390400
transform 1 0 36512 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_318
timestamp 1669390400
transform 1 0 36960 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_321
timestamp 1669390400
transform 1 0 37296 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_385
timestamp 1669390400
transform 1 0 44464 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_389
timestamp 1669390400
transform 1 0 44912 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_392
timestamp 1669390400
transform 1 0 45248 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_456
timestamp 1669390400
transform 1 0 52416 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_460
timestamp 1669390400
transform 1 0 52864 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_463
timestamp 1669390400
transform 1 0 53200 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_527
timestamp 1669390400
transform 1 0 60368 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_531
timestamp 1669390400
transform 1 0 60816 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_534
timestamp 1669390400
transform 1 0 61152 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_598
timestamp 1669390400
transform 1 0 68320 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_602
timestamp 1669390400
transform 1 0 68768 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_605
timestamp 1669390400
transform 1 0 69104 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_669
timestamp 1669390400
transform 1 0 76272 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_673
timestamp 1669390400
transform 1 0 76720 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_676
timestamp 1669390400
transform 1 0 77056 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_740
timestamp 1669390400
transform 1 0 84224 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_744
timestamp 1669390400
transform 1 0 84672 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_747
timestamp 1669390400
transform 1 0 85008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_811
timestamp 1669390400
transform 1 0 92176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_815
timestamp 1669390400
transform 1 0 92624 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_818
timestamp 1669390400
transform 1 0 92960 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_882
timestamp 1669390400
transform 1 0 100128 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_886
timestamp 1669390400
transform 1 0 100576 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_889
timestamp 1669390400
transform 1 0 100912 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_953
timestamp 1669390400
transform 1 0 108080 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_957
timestamp 1669390400
transform 1 0 108528 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_960
timestamp 1669390400
transform 1 0 108864 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_992
timestamp 1669390400
transform 1 0 112448 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1008
timestamp 1669390400
transform 1 0 114240 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_1011
timestamp 1669390400
transform 1 0 114576 0 1 92512
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_1027
timestamp 1669390400
transform 1 0 116368 0 1 92512
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_1031
timestamp 1669390400
transform 1 0 116816 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1039
timestamp 1669390400
transform 1 0 117712 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_1043
timestamp 1669390400
transform 1 0 118160 0 1 92512
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_2
timestamp 1669390400
transform 1 0 1568 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_17
timestamp 1669390400
transform 1 0 3248 0 -1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_115_21
timestamp 1669390400
transform 1 0 3696 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_53
timestamp 1669390400
transform 1 0 7280 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_69
timestamp 1669390400
transform 1 0 9072 0 -1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_73
timestamp 1669390400
transform 1 0 9520 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_137
timestamp 1669390400
transform 1 0 16688 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_141
timestamp 1669390400
transform 1 0 17136 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_144
timestamp 1669390400
transform 1 0 17472 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_208
timestamp 1669390400
transform 1 0 24640 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_212
timestamp 1669390400
transform 1 0 25088 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_215
timestamp 1669390400
transform 1 0 25424 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_279
timestamp 1669390400
transform 1 0 32592 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_283
timestamp 1669390400
transform 1 0 33040 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_286
timestamp 1669390400
transform 1 0 33376 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_350
timestamp 1669390400
transform 1 0 40544 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_354
timestamp 1669390400
transform 1 0 40992 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_115_357
timestamp 1669390400
transform 1 0 41328 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_389
timestamp 1669390400
transform 1 0 44912 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_115_405
timestamp 1669390400
transform 1 0 46704 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_413
timestamp 1669390400
transform 1 0 47600 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_417
timestamp 1669390400
transform 1 0 48048 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_424
timestamp 1669390400
transform 1 0 48832 0 -1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_428
timestamp 1669390400
transform 1 0 49280 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_431
timestamp 1669390400
transform 1 0 49616 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_495
timestamp 1669390400
transform 1 0 56784 0 -1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_499
timestamp 1669390400
transform 1 0 57232 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_563
timestamp 1669390400
transform 1 0 64400 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_567
timestamp 1669390400
transform 1 0 64848 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_570
timestamp 1669390400
transform 1 0 65184 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_634
timestamp 1669390400
transform 1 0 72352 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_638
timestamp 1669390400
transform 1 0 72800 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_641
timestamp 1669390400
transform 1 0 73136 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_705
timestamp 1669390400
transform 1 0 80304 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_709
timestamp 1669390400
transform 1 0 80752 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_712
timestamp 1669390400
transform 1 0 81088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_776
timestamp 1669390400
transform 1 0 88256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_780
timestamp 1669390400
transform 1 0 88704 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_783
timestamp 1669390400
transform 1 0 89040 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_847
timestamp 1669390400
transform 1 0 96208 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_851
timestamp 1669390400
transform 1 0 96656 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_854
timestamp 1669390400
transform 1 0 96992 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_918
timestamp 1669390400
transform 1 0 104160 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_922
timestamp 1669390400
transform 1 0 104608 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_925
timestamp 1669390400
transform 1 0 104944 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_989
timestamp 1669390400
transform 1 0 112112 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_993
timestamp 1669390400
transform 1 0 112560 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_115_996
timestamp 1669390400
transform 1 0 112896 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_1028
timestamp 1669390400
transform 1 0 116480 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1044
timestamp 1669390400
transform 1 0 118272 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_2
timestamp 1669390400
transform 1 0 1568 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_6
timestamp 1669390400
transform 1 0 2016 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_8
timestamp 1669390400
transform 1 0 2240 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_15
timestamp 1669390400
transform 1 0 3024 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_19
timestamp 1669390400
transform 1 0 3472 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_37
timestamp 1669390400
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_101
timestamp 1669390400
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_105
timestamp 1669390400
transform 1 0 13104 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_108
timestamp 1669390400
transform 1 0 13440 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_172
timestamp 1669390400
transform 1 0 20608 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_176
timestamp 1669390400
transform 1 0 21056 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_179
timestamp 1669390400
transform 1 0 21392 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_243
timestamp 1669390400
transform 1 0 28560 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_247
timestamp 1669390400
transform 1 0 29008 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_250
timestamp 1669390400
transform 1 0 29344 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_314
timestamp 1669390400
transform 1 0 36512 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_318
timestamp 1669390400
transform 1 0 36960 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_321
timestamp 1669390400
transform 1 0 37296 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_385
timestamp 1669390400
transform 1 0 44464 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_389
timestamp 1669390400
transform 1 0 44912 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_392
timestamp 1669390400
transform 1 0 45248 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_456
timestamp 1669390400
transform 1 0 52416 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_460
timestamp 1669390400
transform 1 0 52864 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_463
timestamp 1669390400
transform 1 0 53200 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_527
timestamp 1669390400
transform 1 0 60368 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_531
timestamp 1669390400
transform 1 0 60816 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_534
timestamp 1669390400
transform 1 0 61152 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_598
timestamp 1669390400
transform 1 0 68320 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_602
timestamp 1669390400
transform 1 0 68768 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_605
timestamp 1669390400
transform 1 0 69104 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_621
timestamp 1669390400
transform 1 0 70896 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_623
timestamp 1669390400
transform 1 0 71120 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_626
timestamp 1669390400
transform 1 0 71456 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_634
timestamp 1669390400
transform 1 0 72352 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_116_666
timestamp 1669390400
transform 1 0 75936 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_676
timestamp 1669390400
transform 1 0 77056 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_740
timestamp 1669390400
transform 1 0 84224 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_744
timestamp 1669390400
transform 1 0 84672 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_747
timestamp 1669390400
transform 1 0 85008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_811
timestamp 1669390400
transform 1 0 92176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_815
timestamp 1669390400
transform 1 0 92624 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_818
timestamp 1669390400
transform 1 0 92960 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_882
timestamp 1669390400
transform 1 0 100128 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_886
timestamp 1669390400
transform 1 0 100576 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_889
timestamp 1669390400
transform 1 0 100912 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_953
timestamp 1669390400
transform 1 0 108080 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_957
timestamp 1669390400
transform 1 0 108528 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_960
timestamp 1669390400
transform 1 0 108864 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_992
timestamp 1669390400
transform 1 0 112448 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1008
timestamp 1669390400
transform 1 0 114240 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1028
timestamp 1669390400
transform 1 0 116480 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1031
timestamp 1669390400
transform 1 0 116816 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_116_1034
timestamp 1669390400
transform 1 0 117152 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_1042
timestamp 1669390400
transform 1 0 118048 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1044
timestamp 1669390400
transform 1 0 118272 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_2
timestamp 1669390400
transform 1 0 1568 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_117_17
timestamp 1669390400
transform 1 0 3248 0 -1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_117_49
timestamp 1669390400
transform 1 0 6832 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_65
timestamp 1669390400
transform 1 0 8624 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_117_69
timestamp 1669390400
transform 1 0 9072 0 -1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_73
timestamp 1669390400
transform 1 0 9520 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_137
timestamp 1669390400
transform 1 0 16688 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_141
timestamp 1669390400
transform 1 0 17136 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_144
timestamp 1669390400
transform 1 0 17472 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_208
timestamp 1669390400
transform 1 0 24640 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_212
timestamp 1669390400
transform 1 0 25088 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_215
timestamp 1669390400
transform 1 0 25424 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_279
timestamp 1669390400
transform 1 0 32592 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_283
timestamp 1669390400
transform 1 0 33040 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_286
timestamp 1669390400
transform 1 0 33376 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_350
timestamp 1669390400
transform 1 0 40544 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_354
timestamp 1669390400
transform 1 0 40992 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_357
timestamp 1669390400
transform 1 0 41328 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_421
timestamp 1669390400
transform 1 0 48496 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_425
timestamp 1669390400
transform 1 0 48944 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_428
timestamp 1669390400
transform 1 0 49280 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_492
timestamp 1669390400
transform 1 0 56448 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_496
timestamp 1669390400
transform 1 0 56896 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_499
timestamp 1669390400
transform 1 0 57232 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_563
timestamp 1669390400
transform 1 0 64400 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_567
timestamp 1669390400
transform 1 0 64848 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_570
timestamp 1669390400
transform 1 0 65184 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_634
timestamp 1669390400
transform 1 0 72352 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_638
timestamp 1669390400
transform 1 0 72800 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_641
timestamp 1669390400
transform 1 0 73136 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_705
timestamp 1669390400
transform 1 0 80304 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_709
timestamp 1669390400
transform 1 0 80752 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_712
timestamp 1669390400
transform 1 0 81088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_776
timestamp 1669390400
transform 1 0 88256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_780
timestamp 1669390400
transform 1 0 88704 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_783
timestamp 1669390400
transform 1 0 89040 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_847
timestamp 1669390400
transform 1 0 96208 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_851
timestamp 1669390400
transform 1 0 96656 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_854
timestamp 1669390400
transform 1 0 96992 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_918
timestamp 1669390400
transform 1 0 104160 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_922
timestamp 1669390400
transform 1 0 104608 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_925
timestamp 1669390400
transform 1 0 104944 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_989
timestamp 1669390400
transform 1 0 112112 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_993
timestamp 1669390400
transform 1 0 112560 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_117_996
timestamp 1669390400
transform 1 0 112896 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1004
timestamp 1669390400
transform 1 0 113792 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1008
timestamp 1669390400
transform 1 0 114240 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_117_1011
timestamp 1669390400
transform 1 0 114576 0 -1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_117_1027
timestamp 1669390400
transform 1 0 116368 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_117_1043
timestamp 1669390400
transform 1 0 118160 0 -1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_2
timestamp 1669390400
transform 1 0 1568 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_34
timestamp 1669390400
transform 1 0 5152 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_37
timestamp 1669390400
transform 1 0 5488 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_101
timestamp 1669390400
transform 1 0 12656 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_105
timestamp 1669390400
transform 1 0 13104 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_108
timestamp 1669390400
transform 1 0 13440 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_172
timestamp 1669390400
transform 1 0 20608 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_176
timestamp 1669390400
transform 1 0 21056 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_179
timestamp 1669390400
transform 1 0 21392 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_243
timestamp 1669390400
transform 1 0 28560 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_247
timestamp 1669390400
transform 1 0 29008 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_250
timestamp 1669390400
transform 1 0 29344 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_314
timestamp 1669390400
transform 1 0 36512 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_318
timestamp 1669390400
transform 1 0 36960 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_321
timestamp 1669390400
transform 1 0 37296 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_385
timestamp 1669390400
transform 1 0 44464 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_389
timestamp 1669390400
transform 1 0 44912 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_392
timestamp 1669390400
transform 1 0 45248 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_456
timestamp 1669390400
transform 1 0 52416 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_460
timestamp 1669390400
transform 1 0 52864 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_463
timestamp 1669390400
transform 1 0 53200 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_527
timestamp 1669390400
transform 1 0 60368 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_531
timestamp 1669390400
transform 1 0 60816 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_534
timestamp 1669390400
transform 1 0 61152 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_598
timestamp 1669390400
transform 1 0 68320 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_602
timestamp 1669390400
transform 1 0 68768 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_605
timestamp 1669390400
transform 1 0 69104 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_669
timestamp 1669390400
transform 1 0 76272 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_673
timestamp 1669390400
transform 1 0 76720 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_676
timestamp 1669390400
transform 1 0 77056 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_740
timestamp 1669390400
transform 1 0 84224 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_744
timestamp 1669390400
transform 1 0 84672 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_747
timestamp 1669390400
transform 1 0 85008 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_811
timestamp 1669390400
transform 1 0 92176 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_815
timestamp 1669390400
transform 1 0 92624 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_818
timestamp 1669390400
transform 1 0 92960 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_882
timestamp 1669390400
transform 1 0 100128 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_886
timestamp 1669390400
transform 1 0 100576 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_889
timestamp 1669390400
transform 1 0 100912 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_953
timestamp 1669390400
transform 1 0 108080 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_957
timestamp 1669390400
transform 1 0 108528 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_960
timestamp 1669390400
transform 1 0 108864 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1024
timestamp 1669390400
transform 1 0 116032 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1028
timestamp 1669390400
transform 1 0 116480 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_1031
timestamp 1669390400
transform 1 0 116816 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1039
timestamp 1669390400
transform 1 0 117712 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_1043
timestamp 1669390400
transform 1 0 118160 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_2
timestamp 1669390400
transform 1 0 1568 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_5
timestamp 1669390400
transform 1 0 1904 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_69
timestamp 1669390400
transform 1 0 9072 0 -1 97216
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_73
timestamp 1669390400
transform 1 0 9520 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_137
timestamp 1669390400
transform 1 0 16688 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_141
timestamp 1669390400
transform 1 0 17136 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_144
timestamp 1669390400
transform 1 0 17472 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_208
timestamp 1669390400
transform 1 0 24640 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_212
timestamp 1669390400
transform 1 0 25088 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_215
timestamp 1669390400
transform 1 0 25424 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_279
timestamp 1669390400
transform 1 0 32592 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_283
timestamp 1669390400
transform 1 0 33040 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_286
timestamp 1669390400
transform 1 0 33376 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_350
timestamp 1669390400
transform 1 0 40544 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_354
timestamp 1669390400
transform 1 0 40992 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_357
timestamp 1669390400
transform 1 0 41328 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_421
timestamp 1669390400
transform 1 0 48496 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_425
timestamp 1669390400
transform 1 0 48944 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_428
timestamp 1669390400
transform 1 0 49280 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_492
timestamp 1669390400
transform 1 0 56448 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_496
timestamp 1669390400
transform 1 0 56896 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_499
timestamp 1669390400
transform 1 0 57232 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_563
timestamp 1669390400
transform 1 0 64400 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_567
timestamp 1669390400
transform 1 0 64848 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_570
timestamp 1669390400
transform 1 0 65184 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_634
timestamp 1669390400
transform 1 0 72352 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_638
timestamp 1669390400
transform 1 0 72800 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_641
timestamp 1669390400
transform 1 0 73136 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_705
timestamp 1669390400
transform 1 0 80304 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_709
timestamp 1669390400
transform 1 0 80752 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_712
timestamp 1669390400
transform 1 0 81088 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_776
timestamp 1669390400
transform 1 0 88256 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_780
timestamp 1669390400
transform 1 0 88704 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_783
timestamp 1669390400
transform 1 0 89040 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_847
timestamp 1669390400
transform 1 0 96208 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_851
timestamp 1669390400
transform 1 0 96656 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_854
timestamp 1669390400
transform 1 0 96992 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_918
timestamp 1669390400
transform 1 0 104160 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_922
timestamp 1669390400
transform 1 0 104608 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_925
timestamp 1669390400
transform 1 0 104944 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_989
timestamp 1669390400
transform 1 0 112112 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_993
timestamp 1669390400
transform 1 0 112560 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_119_996
timestamp 1669390400
transform 1 0 112896 0 -1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_119_1028
timestamp 1669390400
transform 1 0 116480 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1036
timestamp 1669390400
transform 1 0 117376 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1044
timestamp 1669390400
transform 1 0 118272 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_2
timestamp 1669390400
transform 1 0 1568 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_120_19
timestamp 1669390400
transform 1 0 3472 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_37
timestamp 1669390400
transform 1 0 5488 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_101
timestamp 1669390400
transform 1 0 12656 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_105
timestamp 1669390400
transform 1 0 13104 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_108
timestamp 1669390400
transform 1 0 13440 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_172
timestamp 1669390400
transform 1 0 20608 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_176
timestamp 1669390400
transform 1 0 21056 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_179
timestamp 1669390400
transform 1 0 21392 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_243
timestamp 1669390400
transform 1 0 28560 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_247
timestamp 1669390400
transform 1 0 29008 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_250
timestamp 1669390400
transform 1 0 29344 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_314
timestamp 1669390400
transform 1 0 36512 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_318
timestamp 1669390400
transform 1 0 36960 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_321
timestamp 1669390400
transform 1 0 37296 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_385
timestamp 1669390400
transform 1 0 44464 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_389
timestamp 1669390400
transform 1 0 44912 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_392
timestamp 1669390400
transform 1 0 45248 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_456
timestamp 1669390400
transform 1 0 52416 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_460
timestamp 1669390400
transform 1 0 52864 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_463
timestamp 1669390400
transform 1 0 53200 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_527
timestamp 1669390400
transform 1 0 60368 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_531
timestamp 1669390400
transform 1 0 60816 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_534
timestamp 1669390400
transform 1 0 61152 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_598
timestamp 1669390400
transform 1 0 68320 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_602
timestamp 1669390400
transform 1 0 68768 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_605
timestamp 1669390400
transform 1 0 69104 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_669
timestamp 1669390400
transform 1 0 76272 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_673
timestamp 1669390400
transform 1 0 76720 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_676
timestamp 1669390400
transform 1 0 77056 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_740
timestamp 1669390400
transform 1 0 84224 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_744
timestamp 1669390400
transform 1 0 84672 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_747
timestamp 1669390400
transform 1 0 85008 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_811
timestamp 1669390400
transform 1 0 92176 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_815
timestamp 1669390400
transform 1 0 92624 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_818
timestamp 1669390400
transform 1 0 92960 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_882
timestamp 1669390400
transform 1 0 100128 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_886
timestamp 1669390400
transform 1 0 100576 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_889
timestamp 1669390400
transform 1 0 100912 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_953
timestamp 1669390400
transform 1 0 108080 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_957
timestamp 1669390400
transform 1 0 108528 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_960
timestamp 1669390400
transform 1 0 108864 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1024
timestamp 1669390400
transform 1 0 116032 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1028
timestamp 1669390400
transform 1 0 116480 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_120_1031
timestamp 1669390400
transform 1 0 116816 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1039
timestamp 1669390400
transform 1 0 117712 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_120_1043
timestamp 1669390400
transform 1 0 118160 0 1 97216
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_2
timestamp 1669390400
transform 1 0 1568 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_121_17
timestamp 1669390400
transform 1 0 3248 0 -1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_121_49
timestamp 1669390400
transform 1 0 6832 0 -1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_65
timestamp 1669390400
transform 1 0 8624 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_69
timestamp 1669390400
transform 1 0 9072 0 -1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_73
timestamp 1669390400
transform 1 0 9520 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_137
timestamp 1669390400
transform 1 0 16688 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_141
timestamp 1669390400
transform 1 0 17136 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_144
timestamp 1669390400
transform 1 0 17472 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_208
timestamp 1669390400
transform 1 0 24640 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_212
timestamp 1669390400
transform 1 0 25088 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_215
timestamp 1669390400
transform 1 0 25424 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_279
timestamp 1669390400
transform 1 0 32592 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_283
timestamp 1669390400
transform 1 0 33040 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_286
timestamp 1669390400
transform 1 0 33376 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_350
timestamp 1669390400
transform 1 0 40544 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_354
timestamp 1669390400
transform 1 0 40992 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_357
timestamp 1669390400
transform 1 0 41328 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_421
timestamp 1669390400
transform 1 0 48496 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_425
timestamp 1669390400
transform 1 0 48944 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_428
timestamp 1669390400
transform 1 0 49280 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_492
timestamp 1669390400
transform 1 0 56448 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_496
timestamp 1669390400
transform 1 0 56896 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_499
timestamp 1669390400
transform 1 0 57232 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_563
timestamp 1669390400
transform 1 0 64400 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_567
timestamp 1669390400
transform 1 0 64848 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_570
timestamp 1669390400
transform 1 0 65184 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_634
timestamp 1669390400
transform 1 0 72352 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_638
timestamp 1669390400
transform 1 0 72800 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_641
timestamp 1669390400
transform 1 0 73136 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_705
timestamp 1669390400
transform 1 0 80304 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_709
timestamp 1669390400
transform 1 0 80752 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_712
timestamp 1669390400
transform 1 0 81088 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_776
timestamp 1669390400
transform 1 0 88256 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_780
timestamp 1669390400
transform 1 0 88704 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_783
timestamp 1669390400
transform 1 0 89040 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_847
timestamp 1669390400
transform 1 0 96208 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_851
timestamp 1669390400
transform 1 0 96656 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_854
timestamp 1669390400
transform 1 0 96992 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_918
timestamp 1669390400
transform 1 0 104160 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_922
timestamp 1669390400
transform 1 0 104608 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_925
timestamp 1669390400
transform 1 0 104944 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_989
timestamp 1669390400
transform 1 0 112112 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_993
timestamp 1669390400
transform 1 0 112560 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_121_996
timestamp 1669390400
transform 1 0 112896 0 -1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_121_1028
timestamp 1669390400
transform 1 0 116480 0 -1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1044
timestamp 1669390400
transform 1 0 118272 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_2
timestamp 1669390400
transform 1 0 1568 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_5
timestamp 1669390400
transform 1 0 1904 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_15
timestamp 1669390400
transform 1 0 3024 0 1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_122_19
timestamp 1669390400
transform 1 0 3472 0 1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_37
timestamp 1669390400
transform 1 0 5488 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_101
timestamp 1669390400
transform 1 0 12656 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_105
timestamp 1669390400
transform 1 0 13104 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_108
timestamp 1669390400
transform 1 0 13440 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_172
timestamp 1669390400
transform 1 0 20608 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_176
timestamp 1669390400
transform 1 0 21056 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_179
timestamp 1669390400
transform 1 0 21392 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_243
timestamp 1669390400
transform 1 0 28560 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_247
timestamp 1669390400
transform 1 0 29008 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_250
timestamp 1669390400
transform 1 0 29344 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_314
timestamp 1669390400
transform 1 0 36512 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_318
timestamp 1669390400
transform 1 0 36960 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_321
timestamp 1669390400
transform 1 0 37296 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_327
timestamp 1669390400
transform 1 0 37968 0 1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_337
timestamp 1669390400
transform 1 0 39088 0 1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_122_341
timestamp 1669390400
transform 1 0 39536 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_122_373
timestamp 1669390400
transform 1 0 43120 0 1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_389
timestamp 1669390400
transform 1 0 44912 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_392
timestamp 1669390400
transform 1 0 45248 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_456
timestamp 1669390400
transform 1 0 52416 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_460
timestamp 1669390400
transform 1 0 52864 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_463
timestamp 1669390400
transform 1 0 53200 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_527
timestamp 1669390400
transform 1 0 60368 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_531
timestamp 1669390400
transform 1 0 60816 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_534
timestamp 1669390400
transform 1 0 61152 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_598
timestamp 1669390400
transform 1 0 68320 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_602
timestamp 1669390400
transform 1 0 68768 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_605
timestamp 1669390400
transform 1 0 69104 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_669
timestamp 1669390400
transform 1 0 76272 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_673
timestamp 1669390400
transform 1 0 76720 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_676
timestamp 1669390400
transform 1 0 77056 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_740
timestamp 1669390400
transform 1 0 84224 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_744
timestamp 1669390400
transform 1 0 84672 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_747
timestamp 1669390400
transform 1 0 85008 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_811
timestamp 1669390400
transform 1 0 92176 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_815
timestamp 1669390400
transform 1 0 92624 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_818
timestamp 1669390400
transform 1 0 92960 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_882
timestamp 1669390400
transform 1 0 100128 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_886
timestamp 1669390400
transform 1 0 100576 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_889
timestamp 1669390400
transform 1 0 100912 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_953
timestamp 1669390400
transform 1 0 108080 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_957
timestamp 1669390400
transform 1 0 108528 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_960
timestamp 1669390400
transform 1 0 108864 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1024
timestamp 1669390400
transform 1 0 116032 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1028
timestamp 1669390400
transform 1 0 116480 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_122_1031
timestamp 1669390400
transform 1 0 116816 0 1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1039
timestamp 1669390400
transform 1 0 117712 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_1043
timestamp 1669390400
transform 1 0 118160 0 1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_2
timestamp 1669390400
transform 1 0 1568 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_123_19
timestamp 1669390400
transform 1 0 3472 0 -1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_51
timestamp 1669390400
transform 1 0 7056 0 -1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_67
timestamp 1669390400
transform 1 0 8848 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_73
timestamp 1669390400
transform 1 0 9520 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_137
timestamp 1669390400
transform 1 0 16688 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_141
timestamp 1669390400
transform 1 0 17136 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_144
timestamp 1669390400
transform 1 0 17472 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_208
timestamp 1669390400
transform 1 0 24640 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_212
timestamp 1669390400
transform 1 0 25088 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_215
timestamp 1669390400
transform 1 0 25424 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_279
timestamp 1669390400
transform 1 0 32592 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_283
timestamp 1669390400
transform 1 0 33040 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_286
timestamp 1669390400
transform 1 0 33376 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_350
timestamp 1669390400
transform 1 0 40544 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_354
timestamp 1669390400
transform 1 0 40992 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_357
timestamp 1669390400
transform 1 0 41328 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_421
timestamp 1669390400
transform 1 0 48496 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_425
timestamp 1669390400
transform 1 0 48944 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_428
timestamp 1669390400
transform 1 0 49280 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_492
timestamp 1669390400
transform 1 0 56448 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_496
timestamp 1669390400
transform 1 0 56896 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_499
timestamp 1669390400
transform 1 0 57232 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_563
timestamp 1669390400
transform 1 0 64400 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_567
timestamp 1669390400
transform 1 0 64848 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_570
timestamp 1669390400
transform 1 0 65184 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_634
timestamp 1669390400
transform 1 0 72352 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_638
timestamp 1669390400
transform 1 0 72800 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_641
timestamp 1669390400
transform 1 0 73136 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_705
timestamp 1669390400
transform 1 0 80304 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_709
timestamp 1669390400
transform 1 0 80752 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_712
timestamp 1669390400
transform 1 0 81088 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_776
timestamp 1669390400
transform 1 0 88256 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_780
timestamp 1669390400
transform 1 0 88704 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_783
timestamp 1669390400
transform 1 0 89040 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_847
timestamp 1669390400
transform 1 0 96208 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_851
timestamp 1669390400
transform 1 0 96656 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_854
timestamp 1669390400
transform 1 0 96992 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_918
timestamp 1669390400
transform 1 0 104160 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_922
timestamp 1669390400
transform 1 0 104608 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_925
timestamp 1669390400
transform 1 0 104944 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_989
timestamp 1669390400
transform 1 0 112112 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_993
timestamp 1669390400
transform 1 0 112560 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_123_996
timestamp 1669390400
transform 1 0 112896 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1004
timestamp 1669390400
transform 1 0 113792 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1008
timestamp 1669390400
transform 1 0 114240 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_123_1011
timestamp 1669390400
transform 1 0 114576 0 -1 100352
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_1027
timestamp 1669390400
transform 1 0 116368 0 -1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_123_1043
timestamp 1669390400
transform 1 0 118160 0 -1 100352
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_124_2
timestamp 1669390400
transform 1 0 1568 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_34
timestamp 1669390400
transform 1 0 5152 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_37
timestamp 1669390400
transform 1 0 5488 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_101
timestamp 1669390400
transform 1 0 12656 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_105
timestamp 1669390400
transform 1 0 13104 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_108
timestamp 1669390400
transform 1 0 13440 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_172
timestamp 1669390400
transform 1 0 20608 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_176
timestamp 1669390400
transform 1 0 21056 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_179
timestamp 1669390400
transform 1 0 21392 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_243
timestamp 1669390400
transform 1 0 28560 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_247
timestamp 1669390400
transform 1 0 29008 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_250
timestamp 1669390400
transform 1 0 29344 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_314
timestamp 1669390400
transform 1 0 36512 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_318
timestamp 1669390400
transform 1 0 36960 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_321
timestamp 1669390400
transform 1 0 37296 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_385
timestamp 1669390400
transform 1 0 44464 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_389
timestamp 1669390400
transform 1 0 44912 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_392
timestamp 1669390400
transform 1 0 45248 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_456
timestamp 1669390400
transform 1 0 52416 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_460
timestamp 1669390400
transform 1 0 52864 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_463
timestamp 1669390400
transform 1 0 53200 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_527
timestamp 1669390400
transform 1 0 60368 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_531
timestamp 1669390400
transform 1 0 60816 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_534
timestamp 1669390400
transform 1 0 61152 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_598
timestamp 1669390400
transform 1 0 68320 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_602
timestamp 1669390400
transform 1 0 68768 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_605
timestamp 1669390400
transform 1 0 69104 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_669
timestamp 1669390400
transform 1 0 76272 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_673
timestamp 1669390400
transform 1 0 76720 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_676
timestamp 1669390400
transform 1 0 77056 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_740
timestamp 1669390400
transform 1 0 84224 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_744
timestamp 1669390400
transform 1 0 84672 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_747
timestamp 1669390400
transform 1 0 85008 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_811
timestamp 1669390400
transform 1 0 92176 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_815
timestamp 1669390400
transform 1 0 92624 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_818
timestamp 1669390400
transform 1 0 92960 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_882
timestamp 1669390400
transform 1 0 100128 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_886
timestamp 1669390400
transform 1 0 100576 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_889
timestamp 1669390400
transform 1 0 100912 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_953
timestamp 1669390400
transform 1 0 108080 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_957
timestamp 1669390400
transform 1 0 108528 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_960
timestamp 1669390400
transform 1 0 108864 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1024
timestamp 1669390400
transform 1 0 116032 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1028
timestamp 1669390400
transform 1 0 116480 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_124_1031
timestamp 1669390400
transform 1 0 116816 0 1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1039
timestamp 1669390400
transform 1 0 117712 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_124_1043
timestamp 1669390400
transform 1 0 118160 0 1 100352
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_2
timestamp 1669390400
transform 1 0 1568 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_125_7
timestamp 1669390400
transform 1 0 2128 0 -1 101920
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_125_11
timestamp 1669390400
transform 1 0 2576 0 -1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_125_43
timestamp 1669390400
transform 1 0 6160 0 -1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_125_59
timestamp 1669390400
transform 1 0 7952 0 -1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_67
timestamp 1669390400
transform 1 0 8848 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_73
timestamp 1669390400
transform 1 0 9520 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_137
timestamp 1669390400
transform 1 0 16688 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_141
timestamp 1669390400
transform 1 0 17136 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_144
timestamp 1669390400
transform 1 0 17472 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_208
timestamp 1669390400
transform 1 0 24640 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_212
timestamp 1669390400
transform 1 0 25088 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_215
timestamp 1669390400
transform 1 0 25424 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_279
timestamp 1669390400
transform 1 0 32592 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_283
timestamp 1669390400
transform 1 0 33040 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_286
timestamp 1669390400
transform 1 0 33376 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_350
timestamp 1669390400
transform 1 0 40544 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_354
timestamp 1669390400
transform 1 0 40992 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_357
timestamp 1669390400
transform 1 0 41328 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_421
timestamp 1669390400
transform 1 0 48496 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_425
timestamp 1669390400
transform 1 0 48944 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_428
timestamp 1669390400
transform 1 0 49280 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_492
timestamp 1669390400
transform 1 0 56448 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_496
timestamp 1669390400
transform 1 0 56896 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_499
timestamp 1669390400
transform 1 0 57232 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_563
timestamp 1669390400
transform 1 0 64400 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_567
timestamp 1669390400
transform 1 0 64848 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_570
timestamp 1669390400
transform 1 0 65184 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_634
timestamp 1669390400
transform 1 0 72352 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_638
timestamp 1669390400
transform 1 0 72800 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_641
timestamp 1669390400
transform 1 0 73136 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_705
timestamp 1669390400
transform 1 0 80304 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_709
timestamp 1669390400
transform 1 0 80752 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_712
timestamp 1669390400
transform 1 0 81088 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_776
timestamp 1669390400
transform 1 0 88256 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_780
timestamp 1669390400
transform 1 0 88704 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_783
timestamp 1669390400
transform 1 0 89040 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_847
timestamp 1669390400
transform 1 0 96208 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_851
timestamp 1669390400
transform 1 0 96656 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_854
timestamp 1669390400
transform 1 0 96992 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_918
timestamp 1669390400
transform 1 0 104160 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_922
timestamp 1669390400
transform 1 0 104608 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_925
timestamp 1669390400
transform 1 0 104944 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_989
timestamp 1669390400
transform 1 0 112112 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_993
timestamp 1669390400
transform 1 0 112560 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_125_996
timestamp 1669390400
transform 1 0 112896 0 -1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_125_1028
timestamp 1669390400
transform 1 0 116480 0 -1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1036
timestamp 1669390400
transform 1 0 117376 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1044
timestamp 1669390400
transform 1 0 118272 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_2
timestamp 1669390400
transform 1 0 1568 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_19
timestamp 1669390400
transform 1 0 3472 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_37
timestamp 1669390400
transform 1 0 5488 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_101
timestamp 1669390400
transform 1 0 12656 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_105
timestamp 1669390400
transform 1 0 13104 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_108
timestamp 1669390400
transform 1 0 13440 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_172
timestamp 1669390400
transform 1 0 20608 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_176
timestamp 1669390400
transform 1 0 21056 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_179
timestamp 1669390400
transform 1 0 21392 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_243
timestamp 1669390400
transform 1 0 28560 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_247
timestamp 1669390400
transform 1 0 29008 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_250
timestamp 1669390400
transform 1 0 29344 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_314
timestamp 1669390400
transform 1 0 36512 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_318
timestamp 1669390400
transform 1 0 36960 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_321
timestamp 1669390400
transform 1 0 37296 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_385
timestamp 1669390400
transform 1 0 44464 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_389
timestamp 1669390400
transform 1 0 44912 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_392
timestamp 1669390400
transform 1 0 45248 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_456
timestamp 1669390400
transform 1 0 52416 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_460
timestamp 1669390400
transform 1 0 52864 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_463
timestamp 1669390400
transform 1 0 53200 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_527
timestamp 1669390400
transform 1 0 60368 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_531
timestamp 1669390400
transform 1 0 60816 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_534
timestamp 1669390400
transform 1 0 61152 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_598
timestamp 1669390400
transform 1 0 68320 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_602
timestamp 1669390400
transform 1 0 68768 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_605
timestamp 1669390400
transform 1 0 69104 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_669
timestamp 1669390400
transform 1 0 76272 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_673
timestamp 1669390400
transform 1 0 76720 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_676
timestamp 1669390400
transform 1 0 77056 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_740
timestamp 1669390400
transform 1 0 84224 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_744
timestamp 1669390400
transform 1 0 84672 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_747
timestamp 1669390400
transform 1 0 85008 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_811
timestamp 1669390400
transform 1 0 92176 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_815
timestamp 1669390400
transform 1 0 92624 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_818
timestamp 1669390400
transform 1 0 92960 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_882
timestamp 1669390400
transform 1 0 100128 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_886
timestamp 1669390400
transform 1 0 100576 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_889
timestamp 1669390400
transform 1 0 100912 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_953
timestamp 1669390400
transform 1 0 108080 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_957
timestamp 1669390400
transform 1 0 108528 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_126_960
timestamp 1669390400
transform 1 0 108864 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_992
timestamp 1669390400
transform 1 0 112448 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1008
timestamp 1669390400
transform 1 0 114240 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1028
timestamp 1669390400
transform 1 0 116480 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1031
timestamp 1669390400
transform 1 0 116816 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_126_1034
timestamp 1669390400
transform 1 0 117152 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_126_1042
timestamp 1669390400
transform 1 0 118048 0 1 101920
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1044
timestamp 1669390400
transform 1 0 118272 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_2
timestamp 1669390400
transform 1 0 1568 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_17
timestamp 1669390400
transform 1 0 3248 0 -1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_127_21
timestamp 1669390400
transform 1 0 3696 0 -1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_53
timestamp 1669390400
transform 1 0 7280 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_69
timestamp 1669390400
transform 1 0 9072 0 -1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_73
timestamp 1669390400
transform 1 0 9520 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_137
timestamp 1669390400
transform 1 0 16688 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_141
timestamp 1669390400
transform 1 0 17136 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_144
timestamp 1669390400
transform 1 0 17472 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_208
timestamp 1669390400
transform 1 0 24640 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_212
timestamp 1669390400
transform 1 0 25088 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_215
timestamp 1669390400
transform 1 0 25424 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_279
timestamp 1669390400
transform 1 0 32592 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_283
timestamp 1669390400
transform 1 0 33040 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_286
timestamp 1669390400
transform 1 0 33376 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_350
timestamp 1669390400
transform 1 0 40544 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_354
timestamp 1669390400
transform 1 0 40992 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_357
timestamp 1669390400
transform 1 0 41328 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_127_373
timestamp 1669390400
transform 1 0 43120 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_381
timestamp 1669390400
transform 1 0 44016 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_385
timestamp 1669390400
transform 1 0 44464 0 -1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_393
timestamp 1669390400
transform 1 0 45360 0 -1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_397
timestamp 1669390400
transform 1 0 45808 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_127_413
timestamp 1669390400
transform 1 0 47600 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_421
timestamp 1669390400
transform 1 0 48496 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_425
timestamp 1669390400
transform 1 0 48944 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_428
timestamp 1669390400
transform 1 0 49280 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_492
timestamp 1669390400
transform 1 0 56448 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_496
timestamp 1669390400
transform 1 0 56896 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_499
timestamp 1669390400
transform 1 0 57232 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_563
timestamp 1669390400
transform 1 0 64400 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_567
timestamp 1669390400
transform 1 0 64848 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_570
timestamp 1669390400
transform 1 0 65184 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_634
timestamp 1669390400
transform 1 0 72352 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_638
timestamp 1669390400
transform 1 0 72800 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_641
timestamp 1669390400
transform 1 0 73136 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_705
timestamp 1669390400
transform 1 0 80304 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_709
timestamp 1669390400
transform 1 0 80752 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_712
timestamp 1669390400
transform 1 0 81088 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_776
timestamp 1669390400
transform 1 0 88256 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_780
timestamp 1669390400
transform 1 0 88704 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_783
timestamp 1669390400
transform 1 0 89040 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_847
timestamp 1669390400
transform 1 0 96208 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_851
timestamp 1669390400
transform 1 0 96656 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_854
timestamp 1669390400
transform 1 0 96992 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_918
timestamp 1669390400
transform 1 0 104160 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_922
timestamp 1669390400
transform 1 0 104608 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_925
timestamp 1669390400
transform 1 0 104944 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_989
timestamp 1669390400
transform 1 0 112112 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_993
timestamp 1669390400
transform 1 0 112560 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_127_996
timestamp 1669390400
transform 1 0 112896 0 -1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_1028
timestamp 1669390400
transform 1 0 116480 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1044
timestamp 1669390400
transform 1 0 118272 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_128_2
timestamp 1669390400
transform 1 0 1568 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_34
timestamp 1669390400
transform 1 0 5152 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_37
timestamp 1669390400
transform 1 0 5488 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_101
timestamp 1669390400
transform 1 0 12656 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_105
timestamp 1669390400
transform 1 0 13104 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_108
timestamp 1669390400
transform 1 0 13440 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_172
timestamp 1669390400
transform 1 0 20608 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_176
timestamp 1669390400
transform 1 0 21056 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_179
timestamp 1669390400
transform 1 0 21392 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_243
timestamp 1669390400
transform 1 0 28560 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_247
timestamp 1669390400
transform 1 0 29008 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_250
timestamp 1669390400
transform 1 0 29344 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_314
timestamp 1669390400
transform 1 0 36512 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_318
timestamp 1669390400
transform 1 0 36960 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_321
timestamp 1669390400
transform 1 0 37296 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_385
timestamp 1669390400
transform 1 0 44464 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_389
timestamp 1669390400
transform 1 0 44912 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_392
timestamp 1669390400
transform 1 0 45248 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_456
timestamp 1669390400
transform 1 0 52416 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_460
timestamp 1669390400
transform 1 0 52864 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_463
timestamp 1669390400
transform 1 0 53200 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_527
timestamp 1669390400
transform 1 0 60368 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_531
timestamp 1669390400
transform 1 0 60816 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_534
timestamp 1669390400
transform 1 0 61152 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_598
timestamp 1669390400
transform 1 0 68320 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_602
timestamp 1669390400
transform 1 0 68768 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_605
timestamp 1669390400
transform 1 0 69104 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_669
timestamp 1669390400
transform 1 0 76272 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_673
timestamp 1669390400
transform 1 0 76720 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_676
timestamp 1669390400
transform 1 0 77056 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_740
timestamp 1669390400
transform 1 0 84224 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_744
timestamp 1669390400
transform 1 0 84672 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_747
timestamp 1669390400
transform 1 0 85008 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_811
timestamp 1669390400
transform 1 0 92176 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_815
timestamp 1669390400
transform 1 0 92624 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_818
timestamp 1669390400
transform 1 0 92960 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_882
timestamp 1669390400
transform 1 0 100128 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_886
timestamp 1669390400
transform 1 0 100576 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_889
timestamp 1669390400
transform 1 0 100912 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_953
timestamp 1669390400
transform 1 0 108080 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_957
timestamp 1669390400
transform 1 0 108528 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_960
timestamp 1669390400
transform 1 0 108864 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1024
timestamp 1669390400
transform 1 0 116032 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1028
timestamp 1669390400
transform 1 0 116480 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_128_1031
timestamp 1669390400
transform 1 0 116816 0 1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1039
timestamp 1669390400
transform 1 0 117712 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_128_1043
timestamp 1669390400
transform 1 0 118160 0 1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_2
timestamp 1669390400
transform 1 0 1568 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_129_17
timestamp 1669390400
transform 1 0 3248 0 -1 105056
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_129_21
timestamp 1669390400
transform 1 0 3696 0 -1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_53
timestamp 1669390400
transform 1 0 7280 0 -1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_129_69
timestamp 1669390400
transform 1 0 9072 0 -1 105056
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_73
timestamp 1669390400
transform 1 0 9520 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_137
timestamp 1669390400
transform 1 0 16688 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_141
timestamp 1669390400
transform 1 0 17136 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_144
timestamp 1669390400
transform 1 0 17472 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_208
timestamp 1669390400
transform 1 0 24640 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_212
timestamp 1669390400
transform 1 0 25088 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_215
timestamp 1669390400
transform 1 0 25424 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_279
timestamp 1669390400
transform 1 0 32592 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_283
timestamp 1669390400
transform 1 0 33040 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_286
timestamp 1669390400
transform 1 0 33376 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_350
timestamp 1669390400
transform 1 0 40544 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_354
timestamp 1669390400
transform 1 0 40992 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_357
timestamp 1669390400
transform 1 0 41328 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_421
timestamp 1669390400
transform 1 0 48496 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_425
timestamp 1669390400
transform 1 0 48944 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_428
timestamp 1669390400
transform 1 0 49280 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_492
timestamp 1669390400
transform 1 0 56448 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_496
timestamp 1669390400
transform 1 0 56896 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_499
timestamp 1669390400
transform 1 0 57232 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_563
timestamp 1669390400
transform 1 0 64400 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_567
timestamp 1669390400
transform 1 0 64848 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_570
timestamp 1669390400
transform 1 0 65184 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_634
timestamp 1669390400
transform 1 0 72352 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_638
timestamp 1669390400
transform 1 0 72800 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_641
timestamp 1669390400
transform 1 0 73136 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_705
timestamp 1669390400
transform 1 0 80304 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_709
timestamp 1669390400
transform 1 0 80752 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_712
timestamp 1669390400
transform 1 0 81088 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_776
timestamp 1669390400
transform 1 0 88256 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_780
timestamp 1669390400
transform 1 0 88704 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_783
timestamp 1669390400
transform 1 0 89040 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_847
timestamp 1669390400
transform 1 0 96208 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_851
timestamp 1669390400
transform 1 0 96656 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_854
timestamp 1669390400
transform 1 0 96992 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_918
timestamp 1669390400
transform 1 0 104160 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_922
timestamp 1669390400
transform 1 0 104608 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_925
timestamp 1669390400
transform 1 0 104944 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_989
timestamp 1669390400
transform 1 0 112112 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_993
timestamp 1669390400
transform 1 0 112560 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_996
timestamp 1669390400
transform 1 0 112896 0 -1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1012
timestamp 1669390400
transform 1 0 114688 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_129_1029
timestamp 1669390400
transform 1 0 116592 0 -1 105056
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_129_1033
timestamp 1669390400
transform 1 0 117040 0 -1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1041
timestamp 1669390400
transform 1 0 117936 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_130_2
timestamp 1669390400
transform 1 0 1568 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_34
timestamp 1669390400
transform 1 0 5152 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_37
timestamp 1669390400
transform 1 0 5488 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_101
timestamp 1669390400
transform 1 0 12656 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_105
timestamp 1669390400
transform 1 0 13104 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_108
timestamp 1669390400
transform 1 0 13440 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_172
timestamp 1669390400
transform 1 0 20608 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_176
timestamp 1669390400
transform 1 0 21056 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_179
timestamp 1669390400
transform 1 0 21392 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_243
timestamp 1669390400
transform 1 0 28560 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_247
timestamp 1669390400
transform 1 0 29008 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_250
timestamp 1669390400
transform 1 0 29344 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_314
timestamp 1669390400
transform 1 0 36512 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_318
timestamp 1669390400
transform 1 0 36960 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_321
timestamp 1669390400
transform 1 0 37296 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_385
timestamp 1669390400
transform 1 0 44464 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_389
timestamp 1669390400
transform 1 0 44912 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_392
timestamp 1669390400
transform 1 0 45248 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_456
timestamp 1669390400
transform 1 0 52416 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_460
timestamp 1669390400
transform 1 0 52864 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_463
timestamp 1669390400
transform 1 0 53200 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_527
timestamp 1669390400
transform 1 0 60368 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_531
timestamp 1669390400
transform 1 0 60816 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_534
timestamp 1669390400
transform 1 0 61152 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_598
timestamp 1669390400
transform 1 0 68320 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_602
timestamp 1669390400
transform 1 0 68768 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_605
timestamp 1669390400
transform 1 0 69104 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_669
timestamp 1669390400
transform 1 0 76272 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_673
timestamp 1669390400
transform 1 0 76720 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_676
timestamp 1669390400
transform 1 0 77056 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_740
timestamp 1669390400
transform 1 0 84224 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_744
timestamp 1669390400
transform 1 0 84672 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_747
timestamp 1669390400
transform 1 0 85008 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_811
timestamp 1669390400
transform 1 0 92176 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_815
timestamp 1669390400
transform 1 0 92624 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_818
timestamp 1669390400
transform 1 0 92960 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_882
timestamp 1669390400
transform 1 0 100128 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_886
timestamp 1669390400
transform 1 0 100576 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_889
timestamp 1669390400
transform 1 0 100912 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_953
timestamp 1669390400
transform 1 0 108080 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_957
timestamp 1669390400
transform 1 0 108528 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_960
timestamp 1669390400
transform 1 0 108864 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1024
timestamp 1669390400
transform 1 0 116032 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1028
timestamp 1669390400
transform 1 0 116480 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_130_1031
timestamp 1669390400
transform 1 0 116816 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1039
timestamp 1669390400
transform 1 0 117712 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_130_1043
timestamp 1669390400
transform 1 0 118160 0 1 105056
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_2
timestamp 1669390400
transform 1 0 1568 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_66
timestamp 1669390400
transform 1 0 8736 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_70
timestamp 1669390400
transform 1 0 9184 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_73
timestamp 1669390400
transform 1 0 9520 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_137
timestamp 1669390400
transform 1 0 16688 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_141
timestamp 1669390400
transform 1 0 17136 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_144
timestamp 1669390400
transform 1 0 17472 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_208
timestamp 1669390400
transform 1 0 24640 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_212
timestamp 1669390400
transform 1 0 25088 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_215
timestamp 1669390400
transform 1 0 25424 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_279
timestamp 1669390400
transform 1 0 32592 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_283
timestamp 1669390400
transform 1 0 33040 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_286
timestamp 1669390400
transform 1 0 33376 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_350
timestamp 1669390400
transform 1 0 40544 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_354
timestamp 1669390400
transform 1 0 40992 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_357
timestamp 1669390400
transform 1 0 41328 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_421
timestamp 1669390400
transform 1 0 48496 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_425
timestamp 1669390400
transform 1 0 48944 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_428
timestamp 1669390400
transform 1 0 49280 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_492
timestamp 1669390400
transform 1 0 56448 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_496
timestamp 1669390400
transform 1 0 56896 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_499
timestamp 1669390400
transform 1 0 57232 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_563
timestamp 1669390400
transform 1 0 64400 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_567
timestamp 1669390400
transform 1 0 64848 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_570
timestamp 1669390400
transform 1 0 65184 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_634
timestamp 1669390400
transform 1 0 72352 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_638
timestamp 1669390400
transform 1 0 72800 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_641
timestamp 1669390400
transform 1 0 73136 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_705
timestamp 1669390400
transform 1 0 80304 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_709
timestamp 1669390400
transform 1 0 80752 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_712
timestamp 1669390400
transform 1 0 81088 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_776
timestamp 1669390400
transform 1 0 88256 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_780
timestamp 1669390400
transform 1 0 88704 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_783
timestamp 1669390400
transform 1 0 89040 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_847
timestamp 1669390400
transform 1 0 96208 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_851
timestamp 1669390400
transform 1 0 96656 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_854
timestamp 1669390400
transform 1 0 96992 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_918
timestamp 1669390400
transform 1 0 104160 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_922
timestamp 1669390400
transform 1 0 104608 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_925
timestamp 1669390400
transform 1 0 104944 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_989
timestamp 1669390400
transform 1 0 112112 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_993
timestamp 1669390400
transform 1 0 112560 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_131_996
timestamp 1669390400
transform 1 0 112896 0 -1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1004
timestamp 1669390400
transform 1 0 113792 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1008
timestamp 1669390400
transform 1 0 114240 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_131_1011
timestamp 1669390400
transform 1 0 114576 0 -1 106624
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_131_1027
timestamp 1669390400
transform 1 0 116368 0 -1 106624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_131_1043
timestamp 1669390400
transform 1 0 118160 0 -1 106624
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_132_2
timestamp 1669390400
transform 1 0 1568 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_34
timestamp 1669390400
transform 1 0 5152 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_37
timestamp 1669390400
transform 1 0 5488 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_101
timestamp 1669390400
transform 1 0 12656 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_105
timestamp 1669390400
transform 1 0 13104 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_108
timestamp 1669390400
transform 1 0 13440 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_172
timestamp 1669390400
transform 1 0 20608 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_176
timestamp 1669390400
transform 1 0 21056 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_179
timestamp 1669390400
transform 1 0 21392 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_243
timestamp 1669390400
transform 1 0 28560 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_247
timestamp 1669390400
transform 1 0 29008 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_250
timestamp 1669390400
transform 1 0 29344 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_314
timestamp 1669390400
transform 1 0 36512 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_318
timestamp 1669390400
transform 1 0 36960 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_321
timestamp 1669390400
transform 1 0 37296 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_385
timestamp 1669390400
transform 1 0 44464 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_389
timestamp 1669390400
transform 1 0 44912 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_392
timestamp 1669390400
transform 1 0 45248 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_456
timestamp 1669390400
transform 1 0 52416 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_460
timestamp 1669390400
transform 1 0 52864 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_463
timestamp 1669390400
transform 1 0 53200 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_527
timestamp 1669390400
transform 1 0 60368 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_531
timestamp 1669390400
transform 1 0 60816 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_534
timestamp 1669390400
transform 1 0 61152 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_598
timestamp 1669390400
transform 1 0 68320 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_602
timestamp 1669390400
transform 1 0 68768 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_605
timestamp 1669390400
transform 1 0 69104 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_669
timestamp 1669390400
transform 1 0 76272 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_673
timestamp 1669390400
transform 1 0 76720 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_676
timestamp 1669390400
transform 1 0 77056 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_740
timestamp 1669390400
transform 1 0 84224 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_744
timestamp 1669390400
transform 1 0 84672 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_747
timestamp 1669390400
transform 1 0 85008 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_811
timestamp 1669390400
transform 1 0 92176 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_815
timestamp 1669390400
transform 1 0 92624 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_818
timestamp 1669390400
transform 1 0 92960 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_882
timestamp 1669390400
transform 1 0 100128 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_886
timestamp 1669390400
transform 1 0 100576 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_889
timestamp 1669390400
transform 1 0 100912 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_953
timestamp 1669390400
transform 1 0 108080 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_957
timestamp 1669390400
transform 1 0 108528 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_960
timestamp 1669390400
transform 1 0 108864 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1024
timestamp 1669390400
transform 1 0 116032 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1028
timestamp 1669390400
transform 1 0 116480 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_132_1031
timestamp 1669390400
transform 1 0 116816 0 1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1039
timestamp 1669390400
transform 1 0 117712 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1044
timestamp 1669390400
transform 1 0 118272 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_2
timestamp 1669390400
transform 1 0 1568 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_7
timestamp 1669390400
transform 1 0 2128 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_73
timestamp 1669390400
transform 1 0 9520 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_137
timestamp 1669390400
transform 1 0 16688 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_141
timestamp 1669390400
transform 1 0 17136 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_144
timestamp 1669390400
transform 1 0 17472 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_208
timestamp 1669390400
transform 1 0 24640 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_212
timestamp 1669390400
transform 1 0 25088 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_215
timestamp 1669390400
transform 1 0 25424 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_279
timestamp 1669390400
transform 1 0 32592 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_283
timestamp 1669390400
transform 1 0 33040 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_286
timestamp 1669390400
transform 1 0 33376 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_350
timestamp 1669390400
transform 1 0 40544 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_354
timestamp 1669390400
transform 1 0 40992 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_357
timestamp 1669390400
transform 1 0 41328 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_421
timestamp 1669390400
transform 1 0 48496 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_425
timestamp 1669390400
transform 1 0 48944 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_428
timestamp 1669390400
transform 1 0 49280 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_492
timestamp 1669390400
transform 1 0 56448 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_496
timestamp 1669390400
transform 1 0 56896 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_499
timestamp 1669390400
transform 1 0 57232 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_563
timestamp 1669390400
transform 1 0 64400 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_567
timestamp 1669390400
transform 1 0 64848 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_570
timestamp 1669390400
transform 1 0 65184 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_634
timestamp 1669390400
transform 1 0 72352 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_638
timestamp 1669390400
transform 1 0 72800 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_641
timestamp 1669390400
transform 1 0 73136 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_705
timestamp 1669390400
transform 1 0 80304 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_709
timestamp 1669390400
transform 1 0 80752 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_712
timestamp 1669390400
transform 1 0 81088 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_776
timestamp 1669390400
transform 1 0 88256 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_780
timestamp 1669390400
transform 1 0 88704 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_783
timestamp 1669390400
transform 1 0 89040 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_847
timestamp 1669390400
transform 1 0 96208 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_851
timestamp 1669390400
transform 1 0 96656 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_854
timestamp 1669390400
transform 1 0 96992 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_918
timestamp 1669390400
transform 1 0 104160 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_922
timestamp 1669390400
transform 1 0 104608 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_925
timestamp 1669390400
transform 1 0 104944 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_989
timestamp 1669390400
transform 1 0 112112 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_993
timestamp 1669390400
transform 1 0 112560 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_996
timestamp 1669390400
transform 1 0 112896 0 -1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1012
timestamp 1669390400
transform 1 0 114688 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_1029
timestamp 1669390400
transform 1 0 116592 0 -1 108192
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_133_1033
timestamp 1669390400
transform 1 0 117040 0 -1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1041
timestamp 1669390400
transform 1 0 117936 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_134_2
timestamp 1669390400
transform 1 0 1568 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_34
timestamp 1669390400
transform 1 0 5152 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_37
timestamp 1669390400
transform 1 0 5488 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_101
timestamp 1669390400
transform 1 0 12656 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_105
timestamp 1669390400
transform 1 0 13104 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_108
timestamp 1669390400
transform 1 0 13440 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_172
timestamp 1669390400
transform 1 0 20608 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_176
timestamp 1669390400
transform 1 0 21056 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_179
timestamp 1669390400
transform 1 0 21392 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_243
timestamp 1669390400
transform 1 0 28560 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_247
timestamp 1669390400
transform 1 0 29008 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_250
timestamp 1669390400
transform 1 0 29344 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_314
timestamp 1669390400
transform 1 0 36512 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_318
timestamp 1669390400
transform 1 0 36960 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_321
timestamp 1669390400
transform 1 0 37296 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_385
timestamp 1669390400
transform 1 0 44464 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_389
timestamp 1669390400
transform 1 0 44912 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_392
timestamp 1669390400
transform 1 0 45248 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_456
timestamp 1669390400
transform 1 0 52416 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_460
timestamp 1669390400
transform 1 0 52864 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_463
timestamp 1669390400
transform 1 0 53200 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_527
timestamp 1669390400
transform 1 0 60368 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_531
timestamp 1669390400
transform 1 0 60816 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_534
timestamp 1669390400
transform 1 0 61152 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_598
timestamp 1669390400
transform 1 0 68320 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_602
timestamp 1669390400
transform 1 0 68768 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_605
timestamp 1669390400
transform 1 0 69104 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_669
timestamp 1669390400
transform 1 0 76272 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_673
timestamp 1669390400
transform 1 0 76720 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_676
timestamp 1669390400
transform 1 0 77056 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_740
timestamp 1669390400
transform 1 0 84224 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_744
timestamp 1669390400
transform 1 0 84672 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_747
timestamp 1669390400
transform 1 0 85008 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_811
timestamp 1669390400
transform 1 0 92176 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_815
timestamp 1669390400
transform 1 0 92624 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_818
timestamp 1669390400
transform 1 0 92960 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_882
timestamp 1669390400
transform 1 0 100128 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_886
timestamp 1669390400
transform 1 0 100576 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_889
timestamp 1669390400
transform 1 0 100912 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_953
timestamp 1669390400
transform 1 0 108080 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_957
timestamp 1669390400
transform 1 0 108528 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_960
timestamp 1669390400
transform 1 0 108864 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1024
timestamp 1669390400
transform 1 0 116032 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1028
timestamp 1669390400
transform 1 0 116480 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_134_1031
timestamp 1669390400
transform 1 0 116816 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1039
timestamp 1669390400
transform 1 0 117712 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_134_1043
timestamp 1669390400
transform 1 0 118160 0 1 108192
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_2
timestamp 1669390400
transform 1 0 1568 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_66
timestamp 1669390400
transform 1 0 8736 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_70
timestamp 1669390400
transform 1 0 9184 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_73
timestamp 1669390400
transform 1 0 9520 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_137
timestamp 1669390400
transform 1 0 16688 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_141
timestamp 1669390400
transform 1 0 17136 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_144
timestamp 1669390400
transform 1 0 17472 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_208
timestamp 1669390400
transform 1 0 24640 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_212
timestamp 1669390400
transform 1 0 25088 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_215
timestamp 1669390400
transform 1 0 25424 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_279
timestamp 1669390400
transform 1 0 32592 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_283
timestamp 1669390400
transform 1 0 33040 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_286
timestamp 1669390400
transform 1 0 33376 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_350
timestamp 1669390400
transform 1 0 40544 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_354
timestamp 1669390400
transform 1 0 40992 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_357
timestamp 1669390400
transform 1 0 41328 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_421
timestamp 1669390400
transform 1 0 48496 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_425
timestamp 1669390400
transform 1 0 48944 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_428
timestamp 1669390400
transform 1 0 49280 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_492
timestamp 1669390400
transform 1 0 56448 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_496
timestamp 1669390400
transform 1 0 56896 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_499
timestamp 1669390400
transform 1 0 57232 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_563
timestamp 1669390400
transform 1 0 64400 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_567
timestamp 1669390400
transform 1 0 64848 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_570
timestamp 1669390400
transform 1 0 65184 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_634
timestamp 1669390400
transform 1 0 72352 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_638
timestamp 1669390400
transform 1 0 72800 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_641
timestamp 1669390400
transform 1 0 73136 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_705
timestamp 1669390400
transform 1 0 80304 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_709
timestamp 1669390400
transform 1 0 80752 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_712
timestamp 1669390400
transform 1 0 81088 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_776
timestamp 1669390400
transform 1 0 88256 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_780
timestamp 1669390400
transform 1 0 88704 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_783
timestamp 1669390400
transform 1 0 89040 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_847
timestamp 1669390400
transform 1 0 96208 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_851
timestamp 1669390400
transform 1 0 96656 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_854
timestamp 1669390400
transform 1 0 96992 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_918
timestamp 1669390400
transform 1 0 104160 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_922
timestamp 1669390400
transform 1 0 104608 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_925
timestamp 1669390400
transform 1 0 104944 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_989
timestamp 1669390400
transform 1 0 112112 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_993
timestamp 1669390400
transform 1 0 112560 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_135_996
timestamp 1669390400
transform 1 0 112896 0 -1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1012
timestamp 1669390400
transform 1 0 114688 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_1029
timestamp 1669390400
transform 1 0 116592 0 -1 109760
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_135_1033
timestamp 1669390400
transform 1 0 117040 0 -1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1041
timestamp 1669390400
transform 1 0 117936 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_2
timestamp 1669390400
transform 1 0 1568 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_7
timestamp 1669390400
transform 1 0 2128 0 1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_23
timestamp 1669390400
transform 1 0 3920 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_31
timestamp 1669390400
transform 1 0 4816 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_37
timestamp 1669390400
transform 1 0 5488 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_101
timestamp 1669390400
transform 1 0 12656 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_105
timestamp 1669390400
transform 1 0 13104 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_108
timestamp 1669390400
transform 1 0 13440 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_172
timestamp 1669390400
transform 1 0 20608 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_176
timestamp 1669390400
transform 1 0 21056 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_179
timestamp 1669390400
transform 1 0 21392 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_243
timestamp 1669390400
transform 1 0 28560 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_247
timestamp 1669390400
transform 1 0 29008 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_250
timestamp 1669390400
transform 1 0 29344 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_314
timestamp 1669390400
transform 1 0 36512 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_318
timestamp 1669390400
transform 1 0 36960 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_321
timestamp 1669390400
transform 1 0 37296 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_385
timestamp 1669390400
transform 1 0 44464 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_389
timestamp 1669390400
transform 1 0 44912 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_392
timestamp 1669390400
transform 1 0 45248 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_456
timestamp 1669390400
transform 1 0 52416 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_460
timestamp 1669390400
transform 1 0 52864 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_463
timestamp 1669390400
transform 1 0 53200 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_527
timestamp 1669390400
transform 1 0 60368 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_531
timestamp 1669390400
transform 1 0 60816 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_534
timestamp 1669390400
transform 1 0 61152 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_598
timestamp 1669390400
transform 1 0 68320 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_602
timestamp 1669390400
transform 1 0 68768 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_605
timestamp 1669390400
transform 1 0 69104 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_669
timestamp 1669390400
transform 1 0 76272 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_673
timestamp 1669390400
transform 1 0 76720 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_676
timestamp 1669390400
transform 1 0 77056 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_740
timestamp 1669390400
transform 1 0 84224 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_744
timestamp 1669390400
transform 1 0 84672 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_747
timestamp 1669390400
transform 1 0 85008 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_811
timestamp 1669390400
transform 1 0 92176 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_815
timestamp 1669390400
transform 1 0 92624 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_818
timestamp 1669390400
transform 1 0 92960 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_882
timestamp 1669390400
transform 1 0 100128 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_886
timestamp 1669390400
transform 1 0 100576 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_889
timestamp 1669390400
transform 1 0 100912 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_953
timestamp 1669390400
transform 1 0 108080 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_957
timestamp 1669390400
transform 1 0 108528 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_960
timestamp 1669390400
transform 1 0 108864 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1024
timestamp 1669390400
transform 1 0 116032 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1028
timestamp 1669390400
transform 1 0 116480 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_1031
timestamp 1669390400
transform 1 0 116816 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1039
timestamp 1669390400
transform 1 0 117712 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_136_1043
timestamp 1669390400
transform 1 0 118160 0 1 109760
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_2
timestamp 1669390400
transform 1 0 1568 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_5
timestamp 1669390400
transform 1 0 1904 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_69
timestamp 1669390400
transform 1 0 9072 0 -1 111328
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_73
timestamp 1669390400
transform 1 0 9520 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_137
timestamp 1669390400
transform 1 0 16688 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_141
timestamp 1669390400
transform 1 0 17136 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_144
timestamp 1669390400
transform 1 0 17472 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_208
timestamp 1669390400
transform 1 0 24640 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_212
timestamp 1669390400
transform 1 0 25088 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_215
timestamp 1669390400
transform 1 0 25424 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_279
timestamp 1669390400
transform 1 0 32592 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_283
timestamp 1669390400
transform 1 0 33040 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_286
timestamp 1669390400
transform 1 0 33376 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_350
timestamp 1669390400
transform 1 0 40544 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_354
timestamp 1669390400
transform 1 0 40992 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_357
timestamp 1669390400
transform 1 0 41328 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_421
timestamp 1669390400
transform 1 0 48496 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_425
timestamp 1669390400
transform 1 0 48944 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_428
timestamp 1669390400
transform 1 0 49280 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_492
timestamp 1669390400
transform 1 0 56448 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_496
timestamp 1669390400
transform 1 0 56896 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_499
timestamp 1669390400
transform 1 0 57232 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_563
timestamp 1669390400
transform 1 0 64400 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_567
timestamp 1669390400
transform 1 0 64848 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_570
timestamp 1669390400
transform 1 0 65184 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_634
timestamp 1669390400
transform 1 0 72352 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_638
timestamp 1669390400
transform 1 0 72800 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_641
timestamp 1669390400
transform 1 0 73136 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_705
timestamp 1669390400
transform 1 0 80304 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_709
timestamp 1669390400
transform 1 0 80752 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_712
timestamp 1669390400
transform 1 0 81088 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_776
timestamp 1669390400
transform 1 0 88256 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_780
timestamp 1669390400
transform 1 0 88704 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_783
timestamp 1669390400
transform 1 0 89040 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_847
timestamp 1669390400
transform 1 0 96208 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_851
timestamp 1669390400
transform 1 0 96656 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_854
timestamp 1669390400
transform 1 0 96992 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_918
timestamp 1669390400
transform 1 0 104160 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_922
timestamp 1669390400
transform 1 0 104608 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_925
timestamp 1669390400
transform 1 0 104944 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_989
timestamp 1669390400
transform 1 0 112112 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_993
timestamp 1669390400
transform 1 0 112560 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_137_996
timestamp 1669390400
transform 1 0 112896 0 -1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1012
timestamp 1669390400
transform 1 0 114688 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_1027
timestamp 1669390400
transform 1 0 116368 0 -1 111328
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_137_1031
timestamp 1669390400
transform 1 0 116816 0 -1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1039
timestamp 1669390400
transform 1 0 117712 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_1043
timestamp 1669390400
transform 1 0 118160 0 -1 111328
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_2
timestamp 1669390400
transform 1 0 1568 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_138_19
timestamp 1669390400
transform 1 0 3472 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_37
timestamp 1669390400
transform 1 0 5488 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_101
timestamp 1669390400
transform 1 0 12656 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_105
timestamp 1669390400
transform 1 0 13104 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_108
timestamp 1669390400
transform 1 0 13440 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_172
timestamp 1669390400
transform 1 0 20608 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_176
timestamp 1669390400
transform 1 0 21056 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_179
timestamp 1669390400
transform 1 0 21392 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_243
timestamp 1669390400
transform 1 0 28560 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_247
timestamp 1669390400
transform 1 0 29008 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_250
timestamp 1669390400
transform 1 0 29344 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_314
timestamp 1669390400
transform 1 0 36512 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_318
timestamp 1669390400
transform 1 0 36960 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_321
timestamp 1669390400
transform 1 0 37296 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_385
timestamp 1669390400
transform 1 0 44464 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_389
timestamp 1669390400
transform 1 0 44912 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_392
timestamp 1669390400
transform 1 0 45248 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_456
timestamp 1669390400
transform 1 0 52416 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_460
timestamp 1669390400
transform 1 0 52864 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_463
timestamp 1669390400
transform 1 0 53200 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_527
timestamp 1669390400
transform 1 0 60368 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_531
timestamp 1669390400
transform 1 0 60816 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_534
timestamp 1669390400
transform 1 0 61152 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_598
timestamp 1669390400
transform 1 0 68320 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_602
timestamp 1669390400
transform 1 0 68768 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_605
timestamp 1669390400
transform 1 0 69104 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_669
timestamp 1669390400
transform 1 0 76272 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_673
timestamp 1669390400
transform 1 0 76720 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_676
timestamp 1669390400
transform 1 0 77056 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_740
timestamp 1669390400
transform 1 0 84224 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_744
timestamp 1669390400
transform 1 0 84672 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_747
timestamp 1669390400
transform 1 0 85008 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_811
timestamp 1669390400
transform 1 0 92176 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_815
timestamp 1669390400
transform 1 0 92624 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_818
timestamp 1669390400
transform 1 0 92960 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_882
timestamp 1669390400
transform 1 0 100128 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_886
timestamp 1669390400
transform 1 0 100576 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_889
timestamp 1669390400
transform 1 0 100912 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_953
timestamp 1669390400
transform 1 0 108080 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_957
timestamp 1669390400
transform 1 0 108528 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_960
timestamp 1669390400
transform 1 0 108864 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1024
timestamp 1669390400
transform 1 0 116032 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1028
timestamp 1669390400
transform 1 0 116480 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_1031
timestamp 1669390400
transform 1 0 116816 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1039
timestamp 1669390400
transform 1 0 117712 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1044
timestamp 1669390400
transform 1 0 118272 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_2
timestamp 1669390400
transform 1 0 1568 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_139_17
timestamp 1669390400
transform 1 0 3248 0 -1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_139_49
timestamp 1669390400
transform 1 0 6832 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_65
timestamp 1669390400
transform 1 0 8624 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_139_69
timestamp 1669390400
transform 1 0 9072 0 -1 112896
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_73
timestamp 1669390400
transform 1 0 9520 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_137
timestamp 1669390400
transform 1 0 16688 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_141
timestamp 1669390400
transform 1 0 17136 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_144
timestamp 1669390400
transform 1 0 17472 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_208
timestamp 1669390400
transform 1 0 24640 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_212
timestamp 1669390400
transform 1 0 25088 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_215
timestamp 1669390400
transform 1 0 25424 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_279
timestamp 1669390400
transform 1 0 32592 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_283
timestamp 1669390400
transform 1 0 33040 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_286
timestamp 1669390400
transform 1 0 33376 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_350
timestamp 1669390400
transform 1 0 40544 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_354
timestamp 1669390400
transform 1 0 40992 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_357
timestamp 1669390400
transform 1 0 41328 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_421
timestamp 1669390400
transform 1 0 48496 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_425
timestamp 1669390400
transform 1 0 48944 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_428
timestamp 1669390400
transform 1 0 49280 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_492
timestamp 1669390400
transform 1 0 56448 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_496
timestamp 1669390400
transform 1 0 56896 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_499
timestamp 1669390400
transform 1 0 57232 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_563
timestamp 1669390400
transform 1 0 64400 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_567
timestamp 1669390400
transform 1 0 64848 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_570
timestamp 1669390400
transform 1 0 65184 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_634
timestamp 1669390400
transform 1 0 72352 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_638
timestamp 1669390400
transform 1 0 72800 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_641
timestamp 1669390400
transform 1 0 73136 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_705
timestamp 1669390400
transform 1 0 80304 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_709
timestamp 1669390400
transform 1 0 80752 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_712
timestamp 1669390400
transform 1 0 81088 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_776
timestamp 1669390400
transform 1 0 88256 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_780
timestamp 1669390400
transform 1 0 88704 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_783
timestamp 1669390400
transform 1 0 89040 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_847
timestamp 1669390400
transform 1 0 96208 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_851
timestamp 1669390400
transform 1 0 96656 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_854
timestamp 1669390400
transform 1 0 96992 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_918
timestamp 1669390400
transform 1 0 104160 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_922
timestamp 1669390400
transform 1 0 104608 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_925
timestamp 1669390400
transform 1 0 104944 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_989
timestamp 1669390400
transform 1 0 112112 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_993
timestamp 1669390400
transform 1 0 112560 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_139_996
timestamp 1669390400
transform 1 0 112896 0 -1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_139_1028
timestamp 1669390400
transform 1 0 116480 0 -1 112896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1036
timestamp 1669390400
transform 1 0 117376 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1044
timestamp 1669390400
transform 1 0 118272 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_2
timestamp 1669390400
transform 1 0 1568 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_5
timestamp 1669390400
transform 1 0 1904 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_140_15
timestamp 1669390400
transform 1 0 3024 0 1 112896
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_140_19
timestamp 1669390400
transform 1 0 3472 0 1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_37
timestamp 1669390400
transform 1 0 5488 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_101
timestamp 1669390400
transform 1 0 12656 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_105
timestamp 1669390400
transform 1 0 13104 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_108
timestamp 1669390400
transform 1 0 13440 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_172
timestamp 1669390400
transform 1 0 20608 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_176
timestamp 1669390400
transform 1 0 21056 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_179
timestamp 1669390400
transform 1 0 21392 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_243
timestamp 1669390400
transform 1 0 28560 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_247
timestamp 1669390400
transform 1 0 29008 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_250
timestamp 1669390400
transform 1 0 29344 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_314
timestamp 1669390400
transform 1 0 36512 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_318
timestamp 1669390400
transform 1 0 36960 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_321
timestamp 1669390400
transform 1 0 37296 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_385
timestamp 1669390400
transform 1 0 44464 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_389
timestamp 1669390400
transform 1 0 44912 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_392
timestamp 1669390400
transform 1 0 45248 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_456
timestamp 1669390400
transform 1 0 52416 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_460
timestamp 1669390400
transform 1 0 52864 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_463
timestamp 1669390400
transform 1 0 53200 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_527
timestamp 1669390400
transform 1 0 60368 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_531
timestamp 1669390400
transform 1 0 60816 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_534
timestamp 1669390400
transform 1 0 61152 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_598
timestamp 1669390400
transform 1 0 68320 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_602
timestamp 1669390400
transform 1 0 68768 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_605
timestamp 1669390400
transform 1 0 69104 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_669
timestamp 1669390400
transform 1 0 76272 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_673
timestamp 1669390400
transform 1 0 76720 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_676
timestamp 1669390400
transform 1 0 77056 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_740
timestamp 1669390400
transform 1 0 84224 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_744
timestamp 1669390400
transform 1 0 84672 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_747
timestamp 1669390400
transform 1 0 85008 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_811
timestamp 1669390400
transform 1 0 92176 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_815
timestamp 1669390400
transform 1 0 92624 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_818
timestamp 1669390400
transform 1 0 92960 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_882
timestamp 1669390400
transform 1 0 100128 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_886
timestamp 1669390400
transform 1 0 100576 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_889
timestamp 1669390400
transform 1 0 100912 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_953
timestamp 1669390400
transform 1 0 108080 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_957
timestamp 1669390400
transform 1 0 108528 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_960
timestamp 1669390400
transform 1 0 108864 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1024
timestamp 1669390400
transform 1 0 116032 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1028
timestamp 1669390400
transform 1 0 116480 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_140_1031
timestamp 1669390400
transform 1 0 116816 0 1 112896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1039
timestamp 1669390400
transform 1 0 117712 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_140_1043
timestamp 1669390400
transform 1 0 118160 0 1 112896
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_2
timestamp 1669390400
transform 1 0 1568 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_19
timestamp 1669390400
transform 1 0 3472 0 -1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_141_23
timestamp 1669390400
transform 1 0 3920 0 -1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_141_55
timestamp 1669390400
transform 1 0 7504 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_73
timestamp 1669390400
transform 1 0 9520 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_137
timestamp 1669390400
transform 1 0 16688 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_141
timestamp 1669390400
transform 1 0 17136 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_144
timestamp 1669390400
transform 1 0 17472 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_208
timestamp 1669390400
transform 1 0 24640 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_212
timestamp 1669390400
transform 1 0 25088 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_215
timestamp 1669390400
transform 1 0 25424 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_279
timestamp 1669390400
transform 1 0 32592 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_283
timestamp 1669390400
transform 1 0 33040 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_286
timestamp 1669390400
transform 1 0 33376 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_350
timestamp 1669390400
transform 1 0 40544 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_354
timestamp 1669390400
transform 1 0 40992 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_357
timestamp 1669390400
transform 1 0 41328 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_421
timestamp 1669390400
transform 1 0 48496 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_425
timestamp 1669390400
transform 1 0 48944 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_428
timestamp 1669390400
transform 1 0 49280 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_492
timestamp 1669390400
transform 1 0 56448 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_496
timestamp 1669390400
transform 1 0 56896 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_141_499
timestamp 1669390400
transform 1 0 57232 0 -1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_141_531
timestamp 1669390400
transform 1 0 60816 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_141_547
timestamp 1669390400
transform 1 0 62608 0 -1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_555
timestamp 1669390400
transform 1 0 63504 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_559
timestamp 1669390400
transform 1 0 63952 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_562
timestamp 1669390400
transform 1 0 64288 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_566
timestamp 1669390400
transform 1 0 64736 0 -1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_570
timestamp 1669390400
transform 1 0 65184 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_634
timestamp 1669390400
transform 1 0 72352 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_638
timestamp 1669390400
transform 1 0 72800 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_641
timestamp 1669390400
transform 1 0 73136 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_705
timestamp 1669390400
transform 1 0 80304 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_709
timestamp 1669390400
transform 1 0 80752 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_712
timestamp 1669390400
transform 1 0 81088 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_776
timestamp 1669390400
transform 1 0 88256 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_780
timestamp 1669390400
transform 1 0 88704 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_783
timestamp 1669390400
transform 1 0 89040 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_847
timestamp 1669390400
transform 1 0 96208 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_851
timestamp 1669390400
transform 1 0 96656 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_854
timestamp 1669390400
transform 1 0 96992 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_918
timestamp 1669390400
transform 1 0 104160 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_922
timestamp 1669390400
transform 1 0 104608 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_925
timestamp 1669390400
transform 1 0 104944 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_989
timestamp 1669390400
transform 1 0 112112 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_993
timestamp 1669390400
transform 1 0 112560 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_141_996
timestamp 1669390400
transform 1 0 112896 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1012
timestamp 1669390400
transform 1 0 114688 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_1027
timestamp 1669390400
transform 1 0 116368 0 -1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_1031
timestamp 1669390400
transform 1 0 116816 0 -1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_141_1035
timestamp 1669390400
transform 1 0 117264 0 -1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_1043
timestamp 1669390400
transform 1 0 118160 0 -1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_2
timestamp 1669390400
transform 1 0 1568 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_17
timestamp 1669390400
transform 1 0 3248 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_25
timestamp 1669390400
transform 1 0 4144 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_29
timestamp 1669390400
transform 1 0 4592 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_33
timestamp 1669390400
transform 1 0 5040 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_37
timestamp 1669390400
transform 1 0 5488 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_69
timestamp 1669390400
transform 1 0 9072 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_85
timestamp 1669390400
transform 1 0 10864 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_87
timestamp 1669390400
transform 1 0 11088 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_96
timestamp 1669390400
transform 1 0 12096 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_100
timestamp 1669390400
transform 1 0 12544 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_104
timestamp 1669390400
transform 1 0 12992 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_108
timestamp 1669390400
transform 1 0 13440 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_172
timestamp 1669390400
transform 1 0 20608 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_176
timestamp 1669390400
transform 1 0 21056 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_179
timestamp 1669390400
transform 1 0 21392 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_195
timestamp 1669390400
transform 1 0 23184 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_199
timestamp 1669390400
transform 1 0 23632 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_202
timestamp 1669390400
transform 1 0 23968 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_234
timestamp 1669390400
transform 1 0 27552 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_242
timestamp 1669390400
transform 1 0 28448 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_246
timestamp 1669390400
transform 1 0 28896 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_250
timestamp 1669390400
transform 1 0 29344 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_282
timestamp 1669390400
transform 1 0 32928 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_286
timestamp 1669390400
transform 1 0 33376 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_288
timestamp 1669390400
transform 1 0 33600 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_303
timestamp 1669390400
transform 1 0 35280 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_307
timestamp 1669390400
transform 1 0 35728 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_317
timestamp 1669390400
transform 1 0 36848 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_321
timestamp 1669390400
transform 1 0 37296 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_385
timestamp 1669390400
transform 1 0 44464 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_389
timestamp 1669390400
transform 1 0 44912 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_392
timestamp 1669390400
transform 1 0 45248 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_395
timestamp 1669390400
transform 1 0 45584 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_403
timestamp 1669390400
transform 1 0 46480 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_409
timestamp 1669390400
transform 1 0 47152 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_441
timestamp 1669390400
transform 1 0 50736 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_457
timestamp 1669390400
transform 1 0 52528 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_463
timestamp 1669390400
transform 1 0 53200 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_479
timestamp 1669390400
transform 1 0 54992 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_487
timestamp 1669390400
transform 1 0 55888 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_491
timestamp 1669390400
transform 1 0 56336 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_494
timestamp 1669390400
transform 1 0 56672 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_498
timestamp 1669390400
transform 1 0 57120 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_506
timestamp 1669390400
transform 1 0 58016 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_514
timestamp 1669390400
transform 1 0 58912 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_517
timestamp 1669390400
transform 1 0 59248 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_525
timestamp 1669390400
transform 1 0 60144 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_529
timestamp 1669390400
transform 1 0 60592 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_531
timestamp 1669390400
transform 1 0 60816 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_534
timestamp 1669390400
transform 1 0 61152 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_552
timestamp 1669390400
transform 1 0 63168 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_560
timestamp 1669390400
transform 1 0 64064 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_568
timestamp 1669390400
transform 1 0 64960 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_600
timestamp 1669390400
transform 1 0 68544 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_602
timestamp 1669390400
transform 1 0 68768 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_605
timestamp 1669390400
transform 1 0 69104 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_621
timestamp 1669390400
transform 1 0 70896 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_629
timestamp 1669390400
transform 1 0 71792 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_633
timestamp 1669390400
transform 1 0 72240 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_665
timestamp 1669390400
transform 1 0 75824 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_673
timestamp 1669390400
transform 1 0 76720 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_676
timestamp 1669390400
transform 1 0 77056 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_680
timestamp 1669390400
transform 1 0 77504 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_682
timestamp 1669390400
transform 1 0 77728 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_685
timestamp 1669390400
transform 1 0 78064 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_717
timestamp 1669390400
transform 1 0 81648 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_733
timestamp 1669390400
transform 1 0 83440 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_741
timestamp 1669390400
transform 1 0 84336 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_747
timestamp 1669390400
transform 1 0 85008 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_767
timestamp 1669390400
transform 1 0 87248 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_799
timestamp 1669390400
transform 1 0 90832 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_815
timestamp 1669390400
transform 1 0 92624 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_818
timestamp 1669390400
transform 1 0 92960 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_882
timestamp 1669390400
transform 1 0 100128 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_886
timestamp 1669390400
transform 1 0 100576 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_889
timestamp 1669390400
transform 1 0 100912 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_953
timestamp 1669390400
transform 1 0 108080 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_957
timestamp 1669390400
transform 1 0 108528 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_960
timestamp 1669390400
transform 1 0 108864 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_976
timestamp 1669390400
transform 1 0 110656 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_979
timestamp 1669390400
transform 1 0 110992 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_995
timestamp 1669390400
transform 1 0 112784 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1003
timestamp 1669390400
transform 1 0 113680 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_1007
timestamp 1669390400
transform 1 0 114128 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_1011
timestamp 1669390400
transform 1 0 114576 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_1027
timestamp 1669390400
transform 1 0 116368 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1031
timestamp 1669390400
transform 1 0 116816 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1038
timestamp 1669390400
transform 1 0 117600 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_1042
timestamp 1669390400
transform 1 0 118048 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1044
timestamp 1669390400
transform 1 0 118272 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_2
timestamp 1669390400
transform 1 0 1568 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_17
timestamp 1669390400
transform 1 0 3248 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_33
timestamp 1669390400
transform 1 0 5040 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_37
timestamp 1669390400
transform 1 0 5488 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_41
timestamp 1669390400
transform 1 0 5936 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_57
timestamp 1669390400
transform 1 0 7728 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_65
timestamp 1669390400
transform 1 0 8624 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_69
timestamp 1669390400
transform 1 0 9072 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_73
timestamp 1669390400
transform 1 0 9520 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_77
timestamp 1669390400
transform 1 0 9968 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_85
timestamp 1669390400
transform 1 0 10864 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_101
timestamp 1669390400
transform 1 0 12656 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_119
timestamp 1669390400
transform 1 0 14672 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_135
timestamp 1669390400
transform 1 0 16464 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_139
timestamp 1669390400
transform 1 0 16912 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_141
timestamp 1669390400
transform 1 0 17136 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_144
timestamp 1669390400
transform 1 0 17472 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_176
timestamp 1669390400
transform 1 0 21056 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_184
timestamp 1669390400
transform 1 0 21952 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_188
timestamp 1669390400
transform 1 0 22400 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_192
timestamp 1669390400
transform 1 0 22848 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_200
timestamp 1669390400
transform 1 0 23744 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_210
timestamp 1669390400
transform 1 0 24864 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_212
timestamp 1669390400
transform 1 0 25088 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_215
timestamp 1669390400
transform 1 0 25424 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_231
timestamp 1669390400
transform 1 0 27216 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_239
timestamp 1669390400
transform 1 0 28112 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_245
timestamp 1669390400
transform 1 0 28784 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_263
timestamp 1669390400
transform 1 0 30800 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_267
timestamp 1669390400
transform 1 0 31248 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_283
timestamp 1669390400
transform 1 0 33040 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_286
timestamp 1669390400
transform 1 0 33376 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_289
timestamp 1669390400
transform 1 0 33712 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_297
timestamp 1669390400
transform 1 0 34608 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_315
timestamp 1669390400
transform 1 0 36624 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_335
timestamp 1669390400
transform 1 0 38864 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_353
timestamp 1669390400
transform 1 0 40880 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_357
timestamp 1669390400
transform 1 0 41328 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_365
timestamp 1669390400
transform 1 0 42224 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_389
timestamp 1669390400
transform 1 0 44912 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_407
timestamp 1669390400
transform 1 0 46928 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_423
timestamp 1669390400
transform 1 0 48720 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_425
timestamp 1669390400
transform 1 0 48944 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_428
timestamp 1669390400
transform 1 0 49280 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_444
timestamp 1669390400
transform 1 0 51072 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_449
timestamp 1669390400
transform 1 0 51632 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_481
timestamp 1669390400
transform 1 0 55216 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_496
timestamp 1669390400
transform 1 0 56896 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_499
timestamp 1669390400
transform 1 0 57232 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_515
timestamp 1669390400
transform 1 0 59024 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_531
timestamp 1669390400
transform 1 0 60816 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_561
timestamp 1669390400
transform 1 0 64176 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_565
timestamp 1669390400
transform 1 0 64624 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_567
timestamp 1669390400
transform 1 0 64848 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_570
timestamp 1669390400
transform 1 0 65184 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_578
timestamp 1669390400
transform 1 0 66080 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_582
timestamp 1669390400
transform 1 0 66528 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_590
timestamp 1669390400
transform 1 0 67424 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_598
timestamp 1669390400
transform 1 0 68320 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_606
timestamp 1669390400
transform 1 0 69216 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_612
timestamp 1669390400
transform 1 0 69888 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_616
timestamp 1669390400
transform 1 0 70336 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_626
timestamp 1669390400
transform 1 0 71456 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_630
timestamp 1669390400
transform 1 0 71904 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_638
timestamp 1669390400
transform 1 0 72800 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_641
timestamp 1669390400
transform 1 0 73136 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_657
timestamp 1669390400
transform 1 0 74928 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_665
timestamp 1669390400
transform 1 0 75824 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_671
timestamp 1669390400
transform 1 0 76496 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_687
timestamp 1669390400
transform 1 0 78288 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_705
timestamp 1669390400
transform 1 0 80304 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_709
timestamp 1669390400
transform 1 0 80752 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_712
timestamp 1669390400
transform 1 0 81088 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_716
timestamp 1669390400
transform 1 0 81536 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_719
timestamp 1669390400
transform 1 0 81872 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_737
timestamp 1669390400
transform 1 0 83888 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_741
timestamp 1669390400
transform 1 0 84336 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_751
timestamp 1669390400
transform 1 0 85456 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_755
timestamp 1669390400
transform 1 0 85904 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_771
timestamp 1669390400
transform 1 0 87696 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_775
timestamp 1669390400
transform 1 0 88144 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_779
timestamp 1669390400
transform 1 0 88592 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_783
timestamp 1669390400
transform 1 0 89040 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_847
timestamp 1669390400
transform 1 0 96208 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_851
timestamp 1669390400
transform 1 0 96656 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_854
timestamp 1669390400
transform 1 0 96992 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_870
timestamp 1669390400
transform 1 0 98784 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_878
timestamp 1669390400
transform 1 0 99680 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_882
timestamp 1669390400
transform 1 0 100128 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_884
timestamp 1669390400
transform 1 0 100352 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_887
timestamp 1669390400
transform 1 0 100688 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_903
timestamp 1669390400
transform 1 0 102480 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_919
timestamp 1669390400
transform 1 0 104272 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_925
timestamp 1669390400
transform 1 0 104944 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_959
timestamp 1669390400
transform 1 0 108752 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_977
timestamp 1669390400
transform 1 0 110768 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_993
timestamp 1669390400
transform 1 0 112560 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_996
timestamp 1669390400
transform 1 0 112896 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1012
timestamp 1669390400
transform 1 0 114688 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1027
timestamp 1669390400
transform 1 0 116368 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1043
timestamp 1669390400
transform 1 0 118160 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_2
timestamp 1669390400
transform 1 0 1568 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_19
timestamp 1669390400
transform 1 0 3472 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_27
timestamp 1669390400
transform 1 0 4368 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_33
timestamp 1669390400
transform 1 0 5040 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_37
timestamp 1669390400
transform 1 0 5488 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_41
timestamp 1669390400
transform 1 0 5936 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_59
timestamp 1669390400
transform 1 0 7952 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_67
timestamp 1669390400
transform 1 0 8848 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_69
timestamp 1669390400
transform 1 0 9072 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_72
timestamp 1669390400
transform 1 0 9408 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_74
timestamp 1669390400
transform 1 0 9632 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_77
timestamp 1669390400
transform 1 0 9968 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_95
timestamp 1669390400
transform 1 0 11984 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_99
timestamp 1669390400
transform 1 0 12432 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_103
timestamp 1669390400
transform 1 0 12880 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_107
timestamp 1669390400
transform 1 0 13328 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_139
timestamp 1669390400
transform 1 0 16912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_142
timestamp 1669390400
transform 1 0 17248 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_145
timestamp 1669390400
transform 1 0 17584 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_153
timestamp 1669390400
transform 1 0 18480 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_161
timestamp 1669390400
transform 1 0 19376 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_169
timestamp 1669390400
transform 1 0 20272 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_173
timestamp 1669390400
transform 1 0 20720 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_177
timestamp 1669390400
transform 1 0 21168 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_181
timestamp 1669390400
transform 1 0 21616 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_185
timestamp 1669390400
transform 1 0 22064 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_203
timestamp 1669390400
transform 1 0 24080 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_207
timestamp 1669390400
transform 1 0 24528 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_209
timestamp 1669390400
transform 1 0 24752 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_212
timestamp 1669390400
transform 1 0 25088 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_227
timestamp 1669390400
transform 1 0 26768 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_243
timestamp 1669390400
transform 1 0 28560 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_247
timestamp 1669390400
transform 1 0 29008 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_279
timestamp 1669390400
transform 1 0 32592 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_282
timestamp 1669390400
transform 1 0 32928 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_285
timestamp 1669390400
transform 1 0 33264 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_293
timestamp 1669390400
transform 1 0 34160 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_297
timestamp 1669390400
transform 1 0 34608 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_314
timestamp 1669390400
transform 1 0 36512 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_317
timestamp 1669390400
transform 1 0 36848 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_320
timestamp 1669390400
transform 1 0 37184 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_324
timestamp 1669390400
transform 1 0 37632 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_326
timestamp 1669390400
transform 1 0 37856 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_329
timestamp 1669390400
transform 1 0 38192 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_347
timestamp 1669390400
transform 1 0 40208 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_349
timestamp 1669390400
transform 1 0 40432 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_352
timestamp 1669390400
transform 1 0 40768 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_378
timestamp 1669390400
transform 1 0 43680 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_384
timestamp 1669390400
transform 1 0 44352 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_387
timestamp 1669390400
transform 1 0 44688 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_391
timestamp 1669390400
transform 1 0 45136 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_399
timestamp 1669390400
transform 1 0 46032 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_419
timestamp 1669390400
transform 1 0 48272 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_422
timestamp 1669390400
transform 1 0 48608 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_425
timestamp 1669390400
transform 1 0 48944 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_431
timestamp 1669390400
transform 1 0 49616 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_449
timestamp 1669390400
transform 1 0 51632 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_453
timestamp 1669390400
transform 1 0 52080 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_457
timestamp 1669390400
transform 1 0 52528 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_461
timestamp 1669390400
transform 1 0 52976 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_477
timestamp 1669390400
transform 1 0 54768 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_485
timestamp 1669390400
transform 1 0 55664 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_489
timestamp 1669390400
transform 1 0 56112 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_492
timestamp 1669390400
transform 1 0 56448 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_509
timestamp 1669390400
transform 1 0 58352 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_517
timestamp 1669390400
transform 1 0 59248 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_521
timestamp 1669390400
transform 1 0 59696 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_524
timestamp 1669390400
transform 1 0 60032 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_527
timestamp 1669390400
transform 1 0 60368 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_545
timestamp 1669390400
transform 1 0 62384 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_553
timestamp 1669390400
transform 1 0 63280 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_557
timestamp 1669390400
transform 1 0 63728 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_559
timestamp 1669390400
transform 1 0 63952 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_562
timestamp 1669390400
transform 1 0 64288 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_577
timestamp 1669390400
transform 1 0 65968 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_593
timestamp 1669390400
transform 1 0 67760 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_597
timestamp 1669390400
transform 1 0 68208 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_612
timestamp 1669390400
transform 1 0 69888 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_614
timestamp 1669390400
transform 1 0 70112 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_629
timestamp 1669390400
transform 1 0 71792 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_632
timestamp 1669390400
transform 1 0 72128 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_658
timestamp 1669390400
transform 1 0 75040 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_664
timestamp 1669390400
transform 1 0 75712 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_667
timestamp 1669390400
transform 1 0 76048 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_682
timestamp 1669390400
transform 1 0 77728 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_684
timestamp 1669390400
transform 1 0 77952 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_699
timestamp 1669390400
transform 1 0 79632 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_702
timestamp 1669390400
transform 1 0 79968 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_710
timestamp 1669390400
transform 1 0 80864 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_713
timestamp 1669390400
transform 1 0 81200 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_731
timestamp 1669390400
transform 1 0 83216 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_737
timestamp 1669390400
transform 1 0 83888 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_752
timestamp 1669390400
transform 1 0 85568 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_768
timestamp 1669390400
transform 1 0 87360 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_772
timestamp 1669390400
transform 1 0 87808 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_774
timestamp 1669390400
transform 1 0 88032 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_789
timestamp 1669390400
transform 1 0 89712 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_797
timestamp 1669390400
transform 1 0 90608 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_801
timestamp 1669390400
transform 1 0 91056 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_804
timestamp 1669390400
transform 1 0 91392 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_807
timestamp 1669390400
transform 1 0 91728 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_822
timestamp 1669390400
transform 1 0 93408 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_826
timestamp 1669390400
transform 1 0 93856 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_828
timestamp 1669390400
transform 1 0 94080 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_833
timestamp 1669390400
transform 1 0 94640 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_839
timestamp 1669390400
transform 1 0 95312 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_842
timestamp 1669390400
transform 1 0 95648 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_859
timestamp 1669390400
transform 1 0 97552 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_865
timestamp 1669390400
transform 1 0 98224 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_869
timestamp 1669390400
transform 1 0 98672 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_871
timestamp 1669390400
transform 1 0 98896 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_874
timestamp 1669390400
transform 1 0 99232 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_877
timestamp 1669390400
transform 1 0 99568 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_894
timestamp 1669390400
transform 1 0 101472 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_912
timestamp 1669390400
transform 1 0 103488 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_928
timestamp 1669390400
transform 1 0 105280 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_936
timestamp 1669390400
transform 1 0 106176 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_940
timestamp 1669390400
transform 1 0 106624 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_944
timestamp 1669390400
transform 1 0 107072 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_947
timestamp 1669390400
transform 1 0 107408 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_964
timestamp 1669390400
transform 1 0 109312 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_972
timestamp 1669390400
transform 1 0 110208 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_976
timestamp 1669390400
transform 1 0 110656 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_979
timestamp 1669390400
transform 1 0 110992 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_982
timestamp 1669390400
transform 1 0 111328 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_984
timestamp 1669390400
transform 1 0 111552 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1001
timestamp 1669390400
transform 1 0 113456 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1009
timestamp 1669390400
transform 1 0 114352 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1011
timestamp 1669390400
transform 1 0 114576 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1014
timestamp 1669390400
transform 1 0 114912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1017
timestamp 1669390400
transform 1 0 115248 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1034
timestamp 1669390400
transform 1 0 117152 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1038
timestamp 1669390400
transform 1 0 117600 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1042
timestamp 1669390400
transform 1 0 118048 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1044
timestamp 1669390400
transform 1 0 118272 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 118608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 118608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 118608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 118608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 118608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 118608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 118608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 118608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 118608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 118608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 118608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 118608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 118608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 118608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 118608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 118608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 118608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 118608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 118608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 118608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 118608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 118608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 118608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 118608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 118608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 118608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 118608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 118608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 118608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 118608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 118608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 118608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 118608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 118608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 118608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 118608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 118608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 118608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 118608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 118608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 118608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 118608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 118608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 118608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 118608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 118608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 118608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 118608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 118608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 118608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 118608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 118608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 118608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 118608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 118608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 118608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 118608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 118608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 118608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 118608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 118608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 118608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 118608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 118608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 118608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 118608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 118608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 118608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 118608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 118608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 118608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 118608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 118608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 118608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 118608 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 118608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 118608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 118608 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 118608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 118608 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 118608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 118608 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 118608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 118608 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 118608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 118608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 118608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 118608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 118608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 118608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 118608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 118608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 118608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 118608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_188
timestamp 1669390400
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_189
timestamp 1669390400
transform -1 0 118608 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_190
timestamp 1669390400
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_191
timestamp 1669390400
transform -1 0 118608 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_192
timestamp 1669390400
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_193
timestamp 1669390400
transform -1 0 118608 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_194
timestamp 1669390400
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_195
timestamp 1669390400
transform -1 0 118608 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_196
timestamp 1669390400
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_197
timestamp 1669390400
transform -1 0 118608 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_198
timestamp 1669390400
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_199
timestamp 1669390400
transform -1 0 118608 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_200
timestamp 1669390400
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_201
timestamp 1669390400
transform -1 0 118608 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_202
timestamp 1669390400
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_203
timestamp 1669390400
transform -1 0 118608 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_204
timestamp 1669390400
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_205
timestamp 1669390400
transform -1 0 118608 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_206
timestamp 1669390400
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_207
timestamp 1669390400
transform -1 0 118608 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_208
timestamp 1669390400
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_209
timestamp 1669390400
transform -1 0 118608 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_210
timestamp 1669390400
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_211
timestamp 1669390400
transform -1 0 118608 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_212
timestamp 1669390400
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_213
timestamp 1669390400
transform -1 0 118608 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_214
timestamp 1669390400
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_215
timestamp 1669390400
transform -1 0 118608 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_216
timestamp 1669390400
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_217
timestamp 1669390400
transform -1 0 118608 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_218
timestamp 1669390400
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_219
timestamp 1669390400
transform -1 0 118608 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_220
timestamp 1669390400
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_221
timestamp 1669390400
transform -1 0 118608 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_222
timestamp 1669390400
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_223
timestamp 1669390400
transform -1 0 118608 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_224
timestamp 1669390400
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_225
timestamp 1669390400
transform -1 0 118608 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_226
timestamp 1669390400
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_227
timestamp 1669390400
transform -1 0 118608 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_228
timestamp 1669390400
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_229
timestamp 1669390400
transform -1 0 118608 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_230
timestamp 1669390400
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_231
timestamp 1669390400
transform -1 0 118608 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_232
timestamp 1669390400
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_233
timestamp 1669390400
transform -1 0 118608 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_234
timestamp 1669390400
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_235
timestamp 1669390400
transform -1 0 118608 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_236
timestamp 1669390400
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_237
timestamp 1669390400
transform -1 0 118608 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_238
timestamp 1669390400
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_239
timestamp 1669390400
transform -1 0 118608 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_240
timestamp 1669390400
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_241
timestamp 1669390400
transform -1 0 118608 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_242
timestamp 1669390400
transform 1 0 1344 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_243
timestamp 1669390400
transform -1 0 118608 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_244
timestamp 1669390400
transform 1 0 1344 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_245
timestamp 1669390400
transform -1 0 118608 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_246
timestamp 1669390400
transform 1 0 1344 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_247
timestamp 1669390400
transform -1 0 118608 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_248
timestamp 1669390400
transform 1 0 1344 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_249
timestamp 1669390400
transform -1 0 118608 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_250
timestamp 1669390400
transform 1 0 1344 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_251
timestamp 1669390400
transform -1 0 118608 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_252
timestamp 1669390400
transform 1 0 1344 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_253
timestamp 1669390400
transform -1 0 118608 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_254
timestamp 1669390400
transform 1 0 1344 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_255
timestamp 1669390400
transform -1 0 118608 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_256
timestamp 1669390400
transform 1 0 1344 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_257
timestamp 1669390400
transform -1 0 118608 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_258
timestamp 1669390400
transform 1 0 1344 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_259
timestamp 1669390400
transform -1 0 118608 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_260
timestamp 1669390400
transform 1 0 1344 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_261
timestamp 1669390400
transform -1 0 118608 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_262
timestamp 1669390400
transform 1 0 1344 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_263
timestamp 1669390400
transform -1 0 118608 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_264
timestamp 1669390400
transform 1 0 1344 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_265
timestamp 1669390400
transform -1 0 118608 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_266
timestamp 1669390400
transform 1 0 1344 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_267
timestamp 1669390400
transform -1 0 118608 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_268
timestamp 1669390400
transform 1 0 1344 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_269
timestamp 1669390400
transform -1 0 118608 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_270
timestamp 1669390400
transform 1 0 1344 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_271
timestamp 1669390400
transform -1 0 118608 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_272
timestamp 1669390400
transform 1 0 1344 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_273
timestamp 1669390400
transform -1 0 118608 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_274
timestamp 1669390400
transform 1 0 1344 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_275
timestamp 1669390400
transform -1 0 118608 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_276
timestamp 1669390400
transform 1 0 1344 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_277
timestamp 1669390400
transform -1 0 118608 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_278
timestamp 1669390400
transform 1 0 1344 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_279
timestamp 1669390400
transform -1 0 118608 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_280
timestamp 1669390400
transform 1 0 1344 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_281
timestamp 1669390400
transform -1 0 118608 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_282
timestamp 1669390400
transform 1 0 1344 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_283
timestamp 1669390400
transform -1 0 118608 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_284
timestamp 1669390400
transform 1 0 1344 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_285
timestamp 1669390400
transform -1 0 118608 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_286
timestamp 1669390400
transform 1 0 1344 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_287
timestamp 1669390400
transform -1 0 118608 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_288
timestamp 1669390400
transform 1 0 1344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_289
timestamp 1669390400
transform -1 0 118608 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1669390400
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1669390400
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1669390400
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1669390400
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1669390400
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1669390400
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1669390400
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1669390400
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1669390400
transform 1 0 84784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1669390400
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1669390400
transform 1 0 100688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1669390400
transform 1 0 108640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1669390400
transform 1 0 116592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1669390400
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1669390400
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1669390400
transform 1 0 80864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1669390400
transform 1 0 88816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1669390400
transform 1 0 96768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1669390400
transform 1 0 104720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1669390400
transform 1 0 112672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1669390400
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1669390400
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1669390400
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1669390400
transform 1 0 84784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1669390400
transform 1 0 92736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1669390400
transform 1 0 100688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1669390400
transform 1 0 108640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1669390400
transform 1 0 116592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1669390400
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1669390400
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1669390400
transform 1 0 80864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1669390400
transform 1 0 88816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1669390400
transform 1 0 96768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1669390400
transform 1 0 104720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1669390400
transform 1 0 112672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1669390400
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1669390400
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1669390400
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1669390400
transform 1 0 84784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1669390400
transform 1 0 92736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1669390400
transform 1 0 100688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1669390400
transform 1 0 108640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1669390400
transform 1 0 116592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1669390400
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1669390400
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1669390400
transform 1 0 80864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1669390400
transform 1 0 88816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1669390400
transform 1 0 96768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1669390400
transform 1 0 104720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1669390400
transform 1 0 112672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1669390400
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1669390400
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1669390400
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1669390400
transform 1 0 84784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1669390400
transform 1 0 92736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1669390400
transform 1 0 100688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1669390400
transform 1 0 108640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1669390400
transform 1 0 116592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1669390400
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1669390400
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1669390400
transform 1 0 80864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1669390400
transform 1 0 88816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1669390400
transform 1 0 96768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1669390400
transform 1 0 104720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1669390400
transform 1 0 112672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1669390400
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1669390400
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1669390400
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1669390400
transform 1 0 84784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1669390400
transform 1 0 92736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1669390400
transform 1 0 100688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1669390400
transform 1 0 108640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1669390400
transform 1 0 116592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1669390400
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1669390400
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1669390400
transform 1 0 80864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1669390400
transform 1 0 88816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1669390400
transform 1 0 96768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1669390400
transform 1 0 104720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1669390400
transform 1 0 112672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1669390400
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1669390400
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1669390400
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1669390400
transform 1 0 84784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1669390400
transform 1 0 92736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1669390400
transform 1 0 100688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1669390400
transform 1 0 108640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1669390400
transform 1 0 116592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1669390400
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1669390400
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1669390400
transform 1 0 80864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1669390400
transform 1 0 88816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1669390400
transform 1 0 96768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1669390400
transform 1 0 104720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1669390400
transform 1 0 112672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1669390400
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1669390400
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1669390400
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1669390400
transform 1 0 84784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1669390400
transform 1 0 92736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1669390400
transform 1 0 100688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1100
timestamp 1669390400
transform 1 0 108640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1101
timestamp 1669390400
transform 1 0 116592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1102
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1103
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1104
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1105
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1106
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1107
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1108
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1109
timestamp 1669390400
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1110
timestamp 1669390400
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1111
timestamp 1669390400
transform 1 0 80864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1112
timestamp 1669390400
transform 1 0 88816 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1113
timestamp 1669390400
transform 1 0 96768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1114
timestamp 1669390400
transform 1 0 104720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1115
timestamp 1669390400
transform 1 0 112672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1116
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1117
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1118
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1119
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1120
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1121
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1122
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1123
timestamp 1669390400
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1124
timestamp 1669390400
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1125
timestamp 1669390400
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1126
timestamp 1669390400
transform 1 0 84784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1127
timestamp 1669390400
transform 1 0 92736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1128
timestamp 1669390400
transform 1 0 100688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1129
timestamp 1669390400
transform 1 0 108640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1130
timestamp 1669390400
transform 1 0 116592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1131
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1132
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1133
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1134
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1135
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1136
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1137
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1138
timestamp 1669390400
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1139
timestamp 1669390400
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1140
timestamp 1669390400
transform 1 0 80864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1141
timestamp 1669390400
transform 1 0 88816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1142
timestamp 1669390400
transform 1 0 96768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1143
timestamp 1669390400
transform 1 0 104720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1144
timestamp 1669390400
transform 1 0 112672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1145
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1146
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1147
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1148
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1149
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1150
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1151
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1152
timestamp 1669390400
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1153
timestamp 1669390400
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1154
timestamp 1669390400
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1155
timestamp 1669390400
transform 1 0 84784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1156
timestamp 1669390400
transform 1 0 92736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1157
timestamp 1669390400
transform 1 0 100688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1158
timestamp 1669390400
transform 1 0 108640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1159
timestamp 1669390400
transform 1 0 116592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1160
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1161
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1162
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1163
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1164
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1165
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1166
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1167
timestamp 1669390400
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1168
timestamp 1669390400
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1169
timestamp 1669390400
transform 1 0 80864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1170
timestamp 1669390400
transform 1 0 88816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1171
timestamp 1669390400
transform 1 0 96768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1172
timestamp 1669390400
transform 1 0 104720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1173
timestamp 1669390400
transform 1 0 112672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1174
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1175
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1176
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1177
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1178
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1179
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1180
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1181
timestamp 1669390400
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1182
timestamp 1669390400
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1183
timestamp 1669390400
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1184
timestamp 1669390400
transform 1 0 84784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1185
timestamp 1669390400
transform 1 0 92736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1186
timestamp 1669390400
transform 1 0 100688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1187
timestamp 1669390400
transform 1 0 108640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1188
timestamp 1669390400
transform 1 0 116592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1189
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1190
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1191
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1192
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1193
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1194
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1195
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1196
timestamp 1669390400
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1197
timestamp 1669390400
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1198
timestamp 1669390400
transform 1 0 80864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1199
timestamp 1669390400
transform 1 0 88816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1200
timestamp 1669390400
transform 1 0 96768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1201
timestamp 1669390400
transform 1 0 104720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1202
timestamp 1669390400
transform 1 0 112672 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1203
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1204
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1205
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1206
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1207
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1208
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1209
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1210
timestamp 1669390400
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1211
timestamp 1669390400
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1212
timestamp 1669390400
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1213
timestamp 1669390400
transform 1 0 84784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1214
timestamp 1669390400
transform 1 0 92736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1215
timestamp 1669390400
transform 1 0 100688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1216
timestamp 1669390400
transform 1 0 108640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1217
timestamp 1669390400
transform 1 0 116592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1218
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1219
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1220
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1221
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1222
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1223
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1224
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1225
timestamp 1669390400
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1226
timestamp 1669390400
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1227
timestamp 1669390400
transform 1 0 80864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1228
timestamp 1669390400
transform 1 0 88816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1229
timestamp 1669390400
transform 1 0 96768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1230
timestamp 1669390400
transform 1 0 104720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1231
timestamp 1669390400
transform 1 0 112672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1232
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1233
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1234
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1235
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1236
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1237
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1238
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1239
timestamp 1669390400
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1240
timestamp 1669390400
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1241
timestamp 1669390400
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1242
timestamp 1669390400
transform 1 0 84784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1243
timestamp 1669390400
transform 1 0 92736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1244
timestamp 1669390400
transform 1 0 100688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1245
timestamp 1669390400
transform 1 0 108640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1246
timestamp 1669390400
transform 1 0 116592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1247
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1248
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1249
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1250
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1251
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1252
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1253
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1254
timestamp 1669390400
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1255
timestamp 1669390400
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1256
timestamp 1669390400
transform 1 0 80864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1257
timestamp 1669390400
transform 1 0 88816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1258
timestamp 1669390400
transform 1 0 96768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1259
timestamp 1669390400
transform 1 0 104720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1260
timestamp 1669390400
transform 1 0 112672 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1261
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1262
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1263
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1264
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1265
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1266
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1267
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1268
timestamp 1669390400
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1269
timestamp 1669390400
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1270
timestamp 1669390400
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1271
timestamp 1669390400
transform 1 0 84784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1272
timestamp 1669390400
transform 1 0 92736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1273
timestamp 1669390400
transform 1 0 100688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1274
timestamp 1669390400
transform 1 0 108640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1275
timestamp 1669390400
transform 1 0 116592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1276
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1277
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1278
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1279
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1280
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1281
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1282
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1283
timestamp 1669390400
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1284
timestamp 1669390400
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1285
timestamp 1669390400
transform 1 0 80864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1286
timestamp 1669390400
transform 1 0 88816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1287
timestamp 1669390400
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1288
timestamp 1669390400
transform 1 0 104720 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1289
timestamp 1669390400
transform 1 0 112672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1290
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1291
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1292
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1293
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1294
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1295
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1296
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1297
timestamp 1669390400
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1298
timestamp 1669390400
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1299
timestamp 1669390400
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1300
timestamp 1669390400
transform 1 0 84784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1301
timestamp 1669390400
transform 1 0 92736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1302
timestamp 1669390400
transform 1 0 100688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1303
timestamp 1669390400
transform 1 0 108640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1304
timestamp 1669390400
transform 1 0 116592 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1305
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1306
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1307
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1308
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1309
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1310
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1311
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1312
timestamp 1669390400
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1313
timestamp 1669390400
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1314
timestamp 1669390400
transform 1 0 80864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1315
timestamp 1669390400
transform 1 0 88816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1316
timestamp 1669390400
transform 1 0 96768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1317
timestamp 1669390400
transform 1 0 104720 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1318
timestamp 1669390400
transform 1 0 112672 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1319
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1320
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1321
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1322
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1323
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1324
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1325
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1326
timestamp 1669390400
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1327
timestamp 1669390400
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1328
timestamp 1669390400
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1329
timestamp 1669390400
transform 1 0 84784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1330
timestamp 1669390400
transform 1 0 92736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1331
timestamp 1669390400
transform 1 0 100688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1332
timestamp 1669390400
transform 1 0 108640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1333
timestamp 1669390400
transform 1 0 116592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1334
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1335
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1336
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1337
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1338
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1339
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1340
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1341
timestamp 1669390400
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1342
timestamp 1669390400
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1343
timestamp 1669390400
transform 1 0 80864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1344
timestamp 1669390400
transform 1 0 88816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1345
timestamp 1669390400
transform 1 0 96768 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1346
timestamp 1669390400
transform 1 0 104720 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1347
timestamp 1669390400
transform 1 0 112672 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1348
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1349
timestamp 1669390400
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1350
timestamp 1669390400
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1351
timestamp 1669390400
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1352
timestamp 1669390400
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1353
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1354
timestamp 1669390400
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1355
timestamp 1669390400
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1356
timestamp 1669390400
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1357
timestamp 1669390400
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1358
timestamp 1669390400
transform 1 0 84784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1359
timestamp 1669390400
transform 1 0 92736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1360
timestamp 1669390400
transform 1 0 100688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1361
timestamp 1669390400
transform 1 0 108640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1362
timestamp 1669390400
transform 1 0 116592 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1363
timestamp 1669390400
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1364
timestamp 1669390400
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1365
timestamp 1669390400
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1366
timestamp 1669390400
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1367
timestamp 1669390400
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1368
timestamp 1669390400
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1369
timestamp 1669390400
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1370
timestamp 1669390400
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1371
timestamp 1669390400
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1372
timestamp 1669390400
transform 1 0 80864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1373
timestamp 1669390400
transform 1 0 88816 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1374
timestamp 1669390400
transform 1 0 96768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1375
timestamp 1669390400
transform 1 0 104720 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1376
timestamp 1669390400
transform 1 0 112672 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1377
timestamp 1669390400
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1378
timestamp 1669390400
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1379
timestamp 1669390400
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1380
timestamp 1669390400
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1381
timestamp 1669390400
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1382
timestamp 1669390400
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1383
timestamp 1669390400
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1384
timestamp 1669390400
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1385
timestamp 1669390400
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1386
timestamp 1669390400
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1387
timestamp 1669390400
transform 1 0 84784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1388
timestamp 1669390400
transform 1 0 92736 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1389
timestamp 1669390400
transform 1 0 100688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1390
timestamp 1669390400
transform 1 0 108640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1391
timestamp 1669390400
transform 1 0 116592 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1392
timestamp 1669390400
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1393
timestamp 1669390400
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1394
timestamp 1669390400
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1395
timestamp 1669390400
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1396
timestamp 1669390400
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1397
timestamp 1669390400
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1398
timestamp 1669390400
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1399
timestamp 1669390400
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1400
timestamp 1669390400
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1401
timestamp 1669390400
transform 1 0 80864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1402
timestamp 1669390400
transform 1 0 88816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1403
timestamp 1669390400
transform 1 0 96768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1404
timestamp 1669390400
transform 1 0 104720 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1405
timestamp 1669390400
transform 1 0 112672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1406
timestamp 1669390400
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1407
timestamp 1669390400
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1408
timestamp 1669390400
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1409
timestamp 1669390400
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1410
timestamp 1669390400
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1411
timestamp 1669390400
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1412
timestamp 1669390400
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1413
timestamp 1669390400
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1414
timestamp 1669390400
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1415
timestamp 1669390400
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1416
timestamp 1669390400
transform 1 0 84784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1417
timestamp 1669390400
transform 1 0 92736 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1418
timestamp 1669390400
transform 1 0 100688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1419
timestamp 1669390400
transform 1 0 108640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1420
timestamp 1669390400
transform 1 0 116592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1421
timestamp 1669390400
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1422
timestamp 1669390400
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1423
timestamp 1669390400
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1424
timestamp 1669390400
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1425
timestamp 1669390400
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1426
timestamp 1669390400
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1427
timestamp 1669390400
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1428
timestamp 1669390400
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1429
timestamp 1669390400
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1430
timestamp 1669390400
transform 1 0 80864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1431
timestamp 1669390400
transform 1 0 88816 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1432
timestamp 1669390400
transform 1 0 96768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1433
timestamp 1669390400
transform 1 0 104720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1434
timestamp 1669390400
transform 1 0 112672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1435
timestamp 1669390400
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1436
timestamp 1669390400
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1437
timestamp 1669390400
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1438
timestamp 1669390400
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1439
timestamp 1669390400
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1440
timestamp 1669390400
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1441
timestamp 1669390400
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1442
timestamp 1669390400
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1443
timestamp 1669390400
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1444
timestamp 1669390400
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1445
timestamp 1669390400
transform 1 0 84784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1446
timestamp 1669390400
transform 1 0 92736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1447
timestamp 1669390400
transform 1 0 100688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1448
timestamp 1669390400
transform 1 0 108640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1449
timestamp 1669390400
transform 1 0 116592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1450
timestamp 1669390400
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1451
timestamp 1669390400
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1452
timestamp 1669390400
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1453
timestamp 1669390400
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1454
timestamp 1669390400
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1455
timestamp 1669390400
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1456
timestamp 1669390400
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1457
timestamp 1669390400
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1458
timestamp 1669390400
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1459
timestamp 1669390400
transform 1 0 80864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1460
timestamp 1669390400
transform 1 0 88816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1461
timestamp 1669390400
transform 1 0 96768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1462
timestamp 1669390400
transform 1 0 104720 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1463
timestamp 1669390400
transform 1 0 112672 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1464
timestamp 1669390400
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1465
timestamp 1669390400
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1466
timestamp 1669390400
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1467
timestamp 1669390400
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1468
timestamp 1669390400
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1469
timestamp 1669390400
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1470
timestamp 1669390400
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1471
timestamp 1669390400
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1472
timestamp 1669390400
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1473
timestamp 1669390400
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1474
timestamp 1669390400
transform 1 0 84784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1475
timestamp 1669390400
transform 1 0 92736 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1476
timestamp 1669390400
transform 1 0 100688 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1477
timestamp 1669390400
transform 1 0 108640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1478
timestamp 1669390400
transform 1 0 116592 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1479
timestamp 1669390400
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1480
timestamp 1669390400
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1481
timestamp 1669390400
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1482
timestamp 1669390400
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1483
timestamp 1669390400
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1484
timestamp 1669390400
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1485
timestamp 1669390400
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1486
timestamp 1669390400
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1487
timestamp 1669390400
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1488
timestamp 1669390400
transform 1 0 80864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1489
timestamp 1669390400
transform 1 0 88816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1490
timestamp 1669390400
transform 1 0 96768 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1491
timestamp 1669390400
transform 1 0 104720 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1492
timestamp 1669390400
transform 1 0 112672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1493
timestamp 1669390400
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1494
timestamp 1669390400
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1495
timestamp 1669390400
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1496
timestamp 1669390400
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1497
timestamp 1669390400
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1498
timestamp 1669390400
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1499
timestamp 1669390400
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1500
timestamp 1669390400
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1501
timestamp 1669390400
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1502
timestamp 1669390400
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1503
timestamp 1669390400
transform 1 0 84784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1504
timestamp 1669390400
transform 1 0 92736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1505
timestamp 1669390400
transform 1 0 100688 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1506
timestamp 1669390400
transform 1 0 108640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1507
timestamp 1669390400
transform 1 0 116592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1508
timestamp 1669390400
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1509
timestamp 1669390400
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1510
timestamp 1669390400
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1511
timestamp 1669390400
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1512
timestamp 1669390400
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1513
timestamp 1669390400
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1514
timestamp 1669390400
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1515
timestamp 1669390400
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1516
timestamp 1669390400
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1517
timestamp 1669390400
transform 1 0 80864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1518
timestamp 1669390400
transform 1 0 88816 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1519
timestamp 1669390400
transform 1 0 96768 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1520
timestamp 1669390400
transform 1 0 104720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1521
timestamp 1669390400
transform 1 0 112672 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1522
timestamp 1669390400
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1523
timestamp 1669390400
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1524
timestamp 1669390400
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1525
timestamp 1669390400
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1526
timestamp 1669390400
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1527
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1528
timestamp 1669390400
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1529
timestamp 1669390400
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1530
timestamp 1669390400
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1531
timestamp 1669390400
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1532
timestamp 1669390400
transform 1 0 84784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1533
timestamp 1669390400
transform 1 0 92736 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1534
timestamp 1669390400
transform 1 0 100688 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1535
timestamp 1669390400
transform 1 0 108640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1536
timestamp 1669390400
transform 1 0 116592 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1537
timestamp 1669390400
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1538
timestamp 1669390400
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1539
timestamp 1669390400
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1540
timestamp 1669390400
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1541
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1542
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1543
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1544
timestamp 1669390400
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1545
timestamp 1669390400
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1546
timestamp 1669390400
transform 1 0 80864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1547
timestamp 1669390400
transform 1 0 88816 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1548
timestamp 1669390400
transform 1 0 96768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1549
timestamp 1669390400
transform 1 0 104720 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1550
timestamp 1669390400
transform 1 0 112672 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1551
timestamp 1669390400
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1552
timestamp 1669390400
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1553
timestamp 1669390400
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1554
timestamp 1669390400
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1555
timestamp 1669390400
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1556
timestamp 1669390400
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1557
timestamp 1669390400
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1558
timestamp 1669390400
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1559
timestamp 1669390400
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1560
timestamp 1669390400
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1561
timestamp 1669390400
transform 1 0 84784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1562
timestamp 1669390400
transform 1 0 92736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1563
timestamp 1669390400
transform 1 0 100688 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1564
timestamp 1669390400
transform 1 0 108640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1565
timestamp 1669390400
transform 1 0 116592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1566
timestamp 1669390400
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1567
timestamp 1669390400
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1568
timestamp 1669390400
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1569
timestamp 1669390400
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1570
timestamp 1669390400
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1571
timestamp 1669390400
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1572
timestamp 1669390400
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1573
timestamp 1669390400
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1574
timestamp 1669390400
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1575
timestamp 1669390400
transform 1 0 80864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1576
timestamp 1669390400
transform 1 0 88816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1577
timestamp 1669390400
transform 1 0 96768 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1578
timestamp 1669390400
transform 1 0 104720 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1579
timestamp 1669390400
transform 1 0 112672 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1580
timestamp 1669390400
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1581
timestamp 1669390400
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1582
timestamp 1669390400
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1583
timestamp 1669390400
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1584
timestamp 1669390400
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1585
timestamp 1669390400
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1586
timestamp 1669390400
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1587
timestamp 1669390400
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1588
timestamp 1669390400
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1589
timestamp 1669390400
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1590
timestamp 1669390400
transform 1 0 84784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1591
timestamp 1669390400
transform 1 0 92736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1592
timestamp 1669390400
transform 1 0 100688 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1593
timestamp 1669390400
transform 1 0 108640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1594
timestamp 1669390400
transform 1 0 116592 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1595
timestamp 1669390400
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1596
timestamp 1669390400
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1597
timestamp 1669390400
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1598
timestamp 1669390400
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1599
timestamp 1669390400
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1600
timestamp 1669390400
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1601
timestamp 1669390400
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1602
timestamp 1669390400
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1603
timestamp 1669390400
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1604
timestamp 1669390400
transform 1 0 80864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1605
timestamp 1669390400
transform 1 0 88816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1606
timestamp 1669390400
transform 1 0 96768 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1607
timestamp 1669390400
transform 1 0 104720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1608
timestamp 1669390400
transform 1 0 112672 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1609
timestamp 1669390400
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1610
timestamp 1669390400
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1611
timestamp 1669390400
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1612
timestamp 1669390400
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1613
timestamp 1669390400
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1614
timestamp 1669390400
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1615
timestamp 1669390400
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1616
timestamp 1669390400
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1617
timestamp 1669390400
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1618
timestamp 1669390400
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1619
timestamp 1669390400
transform 1 0 84784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1620
timestamp 1669390400
transform 1 0 92736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1621
timestamp 1669390400
transform 1 0 100688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1622
timestamp 1669390400
transform 1 0 108640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1623
timestamp 1669390400
transform 1 0 116592 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1624
timestamp 1669390400
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1625
timestamp 1669390400
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1626
timestamp 1669390400
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1627
timestamp 1669390400
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1628
timestamp 1669390400
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1629
timestamp 1669390400
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1630
timestamp 1669390400
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1631
timestamp 1669390400
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1632
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1633
timestamp 1669390400
transform 1 0 80864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1634
timestamp 1669390400
transform 1 0 88816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1635
timestamp 1669390400
transform 1 0 96768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1636
timestamp 1669390400
transform 1 0 104720 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1637
timestamp 1669390400
transform 1 0 112672 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1638
timestamp 1669390400
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1639
timestamp 1669390400
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1640
timestamp 1669390400
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1641
timestamp 1669390400
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1642
timestamp 1669390400
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1643
timestamp 1669390400
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1644
timestamp 1669390400
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1645
timestamp 1669390400
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1646
timestamp 1669390400
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1647
timestamp 1669390400
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1648
timestamp 1669390400
transform 1 0 84784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1649
timestamp 1669390400
transform 1 0 92736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1650
timestamp 1669390400
transform 1 0 100688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1651
timestamp 1669390400
transform 1 0 108640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1652
timestamp 1669390400
transform 1 0 116592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1653
timestamp 1669390400
transform 1 0 9296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1654
timestamp 1669390400
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1655
timestamp 1669390400
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1656
timestamp 1669390400
transform 1 0 33152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1657
timestamp 1669390400
transform 1 0 41104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1658
timestamp 1669390400
transform 1 0 49056 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1659
timestamp 1669390400
transform 1 0 57008 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1660
timestamp 1669390400
transform 1 0 64960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1661
timestamp 1669390400
transform 1 0 72912 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1662
timestamp 1669390400
transform 1 0 80864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1663
timestamp 1669390400
transform 1 0 88816 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1664
timestamp 1669390400
transform 1 0 96768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1665
timestamp 1669390400
transform 1 0 104720 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1666
timestamp 1669390400
transform 1 0 112672 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1667
timestamp 1669390400
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1668
timestamp 1669390400
transform 1 0 13216 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1669
timestamp 1669390400
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1670
timestamp 1669390400
transform 1 0 29120 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1671
timestamp 1669390400
transform 1 0 37072 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1672
timestamp 1669390400
transform 1 0 45024 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1673
timestamp 1669390400
transform 1 0 52976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1674
timestamp 1669390400
transform 1 0 60928 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1675
timestamp 1669390400
transform 1 0 68880 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1676
timestamp 1669390400
transform 1 0 76832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1677
timestamp 1669390400
transform 1 0 84784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1678
timestamp 1669390400
transform 1 0 92736 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1679
timestamp 1669390400
transform 1 0 100688 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1680
timestamp 1669390400
transform 1 0 108640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1681
timestamp 1669390400
transform 1 0 116592 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1682
timestamp 1669390400
transform 1 0 9296 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1683
timestamp 1669390400
transform 1 0 17248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1684
timestamp 1669390400
transform 1 0 25200 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1685
timestamp 1669390400
transform 1 0 33152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1686
timestamp 1669390400
transform 1 0 41104 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1687
timestamp 1669390400
transform 1 0 49056 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1688
timestamp 1669390400
transform 1 0 57008 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1689
timestamp 1669390400
transform 1 0 64960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1690
timestamp 1669390400
transform 1 0 72912 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1691
timestamp 1669390400
transform 1 0 80864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1692
timestamp 1669390400
transform 1 0 88816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1693
timestamp 1669390400
transform 1 0 96768 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1694
timestamp 1669390400
transform 1 0 104720 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1695
timestamp 1669390400
transform 1 0 112672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1696
timestamp 1669390400
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1697
timestamp 1669390400
transform 1 0 13216 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1698
timestamp 1669390400
transform 1 0 21168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1699
timestamp 1669390400
transform 1 0 29120 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1700
timestamp 1669390400
transform 1 0 37072 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1701
timestamp 1669390400
transform 1 0 45024 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1702
timestamp 1669390400
transform 1 0 52976 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1703
timestamp 1669390400
transform 1 0 60928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1704
timestamp 1669390400
transform 1 0 68880 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1705
timestamp 1669390400
transform 1 0 76832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1706
timestamp 1669390400
transform 1 0 84784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1707
timestamp 1669390400
transform 1 0 92736 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1708
timestamp 1669390400
transform 1 0 100688 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1709
timestamp 1669390400
transform 1 0 108640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1710
timestamp 1669390400
transform 1 0 116592 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1711
timestamp 1669390400
transform 1 0 9296 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1712
timestamp 1669390400
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1713
timestamp 1669390400
transform 1 0 25200 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1714
timestamp 1669390400
transform 1 0 33152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1715
timestamp 1669390400
transform 1 0 41104 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1716
timestamp 1669390400
transform 1 0 49056 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1717
timestamp 1669390400
transform 1 0 57008 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1718
timestamp 1669390400
transform 1 0 64960 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1719
timestamp 1669390400
transform 1 0 72912 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1720
timestamp 1669390400
transform 1 0 80864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1721
timestamp 1669390400
transform 1 0 88816 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1722
timestamp 1669390400
transform 1 0 96768 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1723
timestamp 1669390400
transform 1 0 104720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1724
timestamp 1669390400
transform 1 0 112672 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1725
timestamp 1669390400
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1726
timestamp 1669390400
transform 1 0 13216 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1727
timestamp 1669390400
transform 1 0 21168 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1728
timestamp 1669390400
transform 1 0 29120 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1729
timestamp 1669390400
transform 1 0 37072 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1730
timestamp 1669390400
transform 1 0 45024 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1731
timestamp 1669390400
transform 1 0 52976 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1732
timestamp 1669390400
transform 1 0 60928 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1733
timestamp 1669390400
transform 1 0 68880 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1734
timestamp 1669390400
transform 1 0 76832 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1735
timestamp 1669390400
transform 1 0 84784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1736
timestamp 1669390400
transform 1 0 92736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1737
timestamp 1669390400
transform 1 0 100688 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1738
timestamp 1669390400
transform 1 0 108640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1739
timestamp 1669390400
transform 1 0 116592 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1740
timestamp 1669390400
transform 1 0 9296 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1741
timestamp 1669390400
transform 1 0 17248 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1742
timestamp 1669390400
transform 1 0 25200 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1743
timestamp 1669390400
transform 1 0 33152 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1744
timestamp 1669390400
transform 1 0 41104 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1745
timestamp 1669390400
transform 1 0 49056 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1746
timestamp 1669390400
transform 1 0 57008 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1747
timestamp 1669390400
transform 1 0 64960 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1748
timestamp 1669390400
transform 1 0 72912 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1749
timestamp 1669390400
transform 1 0 80864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1750
timestamp 1669390400
transform 1 0 88816 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1751
timestamp 1669390400
transform 1 0 96768 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1752
timestamp 1669390400
transform 1 0 104720 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1753
timestamp 1669390400
transform 1 0 112672 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1754
timestamp 1669390400
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1755
timestamp 1669390400
transform 1 0 13216 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1756
timestamp 1669390400
transform 1 0 21168 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1757
timestamp 1669390400
transform 1 0 29120 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1758
timestamp 1669390400
transform 1 0 37072 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1759
timestamp 1669390400
transform 1 0 45024 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1760
timestamp 1669390400
transform 1 0 52976 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1761
timestamp 1669390400
transform 1 0 60928 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1762
timestamp 1669390400
transform 1 0 68880 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1763
timestamp 1669390400
transform 1 0 76832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1764
timestamp 1669390400
transform 1 0 84784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1765
timestamp 1669390400
transform 1 0 92736 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1766
timestamp 1669390400
transform 1 0 100688 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1767
timestamp 1669390400
transform 1 0 108640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1768
timestamp 1669390400
transform 1 0 116592 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1769
timestamp 1669390400
transform 1 0 9296 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1770
timestamp 1669390400
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1771
timestamp 1669390400
transform 1 0 25200 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1772
timestamp 1669390400
transform 1 0 33152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1773
timestamp 1669390400
transform 1 0 41104 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1774
timestamp 1669390400
transform 1 0 49056 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1775
timestamp 1669390400
transform 1 0 57008 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1776
timestamp 1669390400
transform 1 0 64960 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1777
timestamp 1669390400
transform 1 0 72912 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1778
timestamp 1669390400
transform 1 0 80864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1779
timestamp 1669390400
transform 1 0 88816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1780
timestamp 1669390400
transform 1 0 96768 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1781
timestamp 1669390400
transform 1 0 104720 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1782
timestamp 1669390400
transform 1 0 112672 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1783
timestamp 1669390400
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1784
timestamp 1669390400
transform 1 0 13216 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1785
timestamp 1669390400
transform 1 0 21168 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1786
timestamp 1669390400
transform 1 0 29120 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1787
timestamp 1669390400
transform 1 0 37072 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1788
timestamp 1669390400
transform 1 0 45024 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1789
timestamp 1669390400
transform 1 0 52976 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1790
timestamp 1669390400
transform 1 0 60928 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1791
timestamp 1669390400
transform 1 0 68880 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1792
timestamp 1669390400
transform 1 0 76832 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1793
timestamp 1669390400
transform 1 0 84784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1794
timestamp 1669390400
transform 1 0 92736 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1795
timestamp 1669390400
transform 1 0 100688 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1796
timestamp 1669390400
transform 1 0 108640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1797
timestamp 1669390400
transform 1 0 116592 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1798
timestamp 1669390400
transform 1 0 9296 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1799
timestamp 1669390400
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1800
timestamp 1669390400
transform 1 0 25200 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1801
timestamp 1669390400
transform 1 0 33152 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1802
timestamp 1669390400
transform 1 0 41104 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1803
timestamp 1669390400
transform 1 0 49056 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1804
timestamp 1669390400
transform 1 0 57008 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1805
timestamp 1669390400
transform 1 0 64960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1806
timestamp 1669390400
transform 1 0 72912 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1807
timestamp 1669390400
transform 1 0 80864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1808
timestamp 1669390400
transform 1 0 88816 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1809
timestamp 1669390400
transform 1 0 96768 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1810
timestamp 1669390400
transform 1 0 104720 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1811
timestamp 1669390400
transform 1 0 112672 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1812
timestamp 1669390400
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1813
timestamp 1669390400
transform 1 0 13216 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1814
timestamp 1669390400
transform 1 0 21168 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1815
timestamp 1669390400
transform 1 0 29120 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1816
timestamp 1669390400
transform 1 0 37072 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1817
timestamp 1669390400
transform 1 0 45024 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1818
timestamp 1669390400
transform 1 0 52976 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1819
timestamp 1669390400
transform 1 0 60928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1820
timestamp 1669390400
transform 1 0 68880 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1821
timestamp 1669390400
transform 1 0 76832 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1822
timestamp 1669390400
transform 1 0 84784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1823
timestamp 1669390400
transform 1 0 92736 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1824
timestamp 1669390400
transform 1 0 100688 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1825
timestamp 1669390400
transform 1 0 108640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1826
timestamp 1669390400
transform 1 0 116592 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1827
timestamp 1669390400
transform 1 0 9296 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1828
timestamp 1669390400
transform 1 0 17248 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1829
timestamp 1669390400
transform 1 0 25200 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1830
timestamp 1669390400
transform 1 0 33152 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1831
timestamp 1669390400
transform 1 0 41104 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1832
timestamp 1669390400
transform 1 0 49056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1833
timestamp 1669390400
transform 1 0 57008 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1834
timestamp 1669390400
transform 1 0 64960 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1835
timestamp 1669390400
transform 1 0 72912 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1836
timestamp 1669390400
transform 1 0 80864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1837
timestamp 1669390400
transform 1 0 88816 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1838
timestamp 1669390400
transform 1 0 96768 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1839
timestamp 1669390400
transform 1 0 104720 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1840
timestamp 1669390400
transform 1 0 112672 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1841
timestamp 1669390400
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1842
timestamp 1669390400
transform 1 0 13216 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1843
timestamp 1669390400
transform 1 0 21168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1844
timestamp 1669390400
transform 1 0 29120 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1845
timestamp 1669390400
transform 1 0 37072 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1846
timestamp 1669390400
transform 1 0 45024 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1847
timestamp 1669390400
transform 1 0 52976 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1848
timestamp 1669390400
transform 1 0 60928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1849
timestamp 1669390400
transform 1 0 68880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1850
timestamp 1669390400
transform 1 0 76832 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1851
timestamp 1669390400
transform 1 0 84784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1852
timestamp 1669390400
transform 1 0 92736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1853
timestamp 1669390400
transform 1 0 100688 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1854
timestamp 1669390400
transform 1 0 108640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1855
timestamp 1669390400
transform 1 0 116592 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1856
timestamp 1669390400
transform 1 0 9296 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1857
timestamp 1669390400
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1858
timestamp 1669390400
transform 1 0 25200 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1859
timestamp 1669390400
transform 1 0 33152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1860
timestamp 1669390400
transform 1 0 41104 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1861
timestamp 1669390400
transform 1 0 49056 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1862
timestamp 1669390400
transform 1 0 57008 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1863
timestamp 1669390400
transform 1 0 64960 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1864
timestamp 1669390400
transform 1 0 72912 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1865
timestamp 1669390400
transform 1 0 80864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1866
timestamp 1669390400
transform 1 0 88816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1867
timestamp 1669390400
transform 1 0 96768 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1868
timestamp 1669390400
transform 1 0 104720 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1869
timestamp 1669390400
transform 1 0 112672 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1870
timestamp 1669390400
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1871
timestamp 1669390400
transform 1 0 13216 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1872
timestamp 1669390400
transform 1 0 21168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1873
timestamp 1669390400
transform 1 0 29120 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1874
timestamp 1669390400
transform 1 0 37072 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1875
timestamp 1669390400
transform 1 0 45024 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1876
timestamp 1669390400
transform 1 0 52976 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1877
timestamp 1669390400
transform 1 0 60928 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1878
timestamp 1669390400
transform 1 0 68880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1879
timestamp 1669390400
transform 1 0 76832 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1880
timestamp 1669390400
transform 1 0 84784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1881
timestamp 1669390400
transform 1 0 92736 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1882
timestamp 1669390400
transform 1 0 100688 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1883
timestamp 1669390400
transform 1 0 108640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1884
timestamp 1669390400
transform 1 0 116592 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1885
timestamp 1669390400
transform 1 0 9296 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1886
timestamp 1669390400
transform 1 0 17248 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1887
timestamp 1669390400
transform 1 0 25200 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1888
timestamp 1669390400
transform 1 0 33152 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1889
timestamp 1669390400
transform 1 0 41104 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1890
timestamp 1669390400
transform 1 0 49056 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1891
timestamp 1669390400
transform 1 0 57008 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1892
timestamp 1669390400
transform 1 0 64960 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1893
timestamp 1669390400
transform 1 0 72912 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1894
timestamp 1669390400
transform 1 0 80864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1895
timestamp 1669390400
transform 1 0 88816 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1896
timestamp 1669390400
transform 1 0 96768 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1897
timestamp 1669390400
transform 1 0 104720 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1898
timestamp 1669390400
transform 1 0 112672 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1899
timestamp 1669390400
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1900
timestamp 1669390400
transform 1 0 13216 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1901
timestamp 1669390400
transform 1 0 21168 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1902
timestamp 1669390400
transform 1 0 29120 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1903
timestamp 1669390400
transform 1 0 37072 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1904
timestamp 1669390400
transform 1 0 45024 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1905
timestamp 1669390400
transform 1 0 52976 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1906
timestamp 1669390400
transform 1 0 60928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1907
timestamp 1669390400
transform 1 0 68880 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1908
timestamp 1669390400
transform 1 0 76832 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1909
timestamp 1669390400
transform 1 0 84784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1910
timestamp 1669390400
transform 1 0 92736 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1911
timestamp 1669390400
transform 1 0 100688 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1912
timestamp 1669390400
transform 1 0 108640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1913
timestamp 1669390400
transform 1 0 116592 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1914
timestamp 1669390400
transform 1 0 9296 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1915
timestamp 1669390400
transform 1 0 17248 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1916
timestamp 1669390400
transform 1 0 25200 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1917
timestamp 1669390400
transform 1 0 33152 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1918
timestamp 1669390400
transform 1 0 41104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1919
timestamp 1669390400
transform 1 0 49056 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1920
timestamp 1669390400
transform 1 0 57008 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1921
timestamp 1669390400
transform 1 0 64960 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1922
timestamp 1669390400
transform 1 0 72912 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1923
timestamp 1669390400
transform 1 0 80864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1924
timestamp 1669390400
transform 1 0 88816 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1925
timestamp 1669390400
transform 1 0 96768 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1926
timestamp 1669390400
transform 1 0 104720 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1927
timestamp 1669390400
transform 1 0 112672 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1928
timestamp 1669390400
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1929
timestamp 1669390400
transform 1 0 13216 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1930
timestamp 1669390400
transform 1 0 21168 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1931
timestamp 1669390400
transform 1 0 29120 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1932
timestamp 1669390400
transform 1 0 37072 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1933
timestamp 1669390400
transform 1 0 45024 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1934
timestamp 1669390400
transform 1 0 52976 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1935
timestamp 1669390400
transform 1 0 60928 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1936
timestamp 1669390400
transform 1 0 68880 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1937
timestamp 1669390400
transform 1 0 76832 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1938
timestamp 1669390400
transform 1 0 84784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1939
timestamp 1669390400
transform 1 0 92736 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1940
timestamp 1669390400
transform 1 0 100688 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1941
timestamp 1669390400
transform 1 0 108640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1942
timestamp 1669390400
transform 1 0 116592 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1943
timestamp 1669390400
transform 1 0 9296 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1944
timestamp 1669390400
transform 1 0 17248 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1945
timestamp 1669390400
transform 1 0 25200 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1946
timestamp 1669390400
transform 1 0 33152 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1947
timestamp 1669390400
transform 1 0 41104 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1948
timestamp 1669390400
transform 1 0 49056 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1949
timestamp 1669390400
transform 1 0 57008 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1950
timestamp 1669390400
transform 1 0 64960 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1951
timestamp 1669390400
transform 1 0 72912 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1952
timestamp 1669390400
transform 1 0 80864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1953
timestamp 1669390400
transform 1 0 88816 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1954
timestamp 1669390400
transform 1 0 96768 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1955
timestamp 1669390400
transform 1 0 104720 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1956
timestamp 1669390400
transform 1 0 112672 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1957
timestamp 1669390400
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1958
timestamp 1669390400
transform 1 0 13216 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1959
timestamp 1669390400
transform 1 0 21168 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1960
timestamp 1669390400
transform 1 0 29120 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1961
timestamp 1669390400
transform 1 0 37072 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1962
timestamp 1669390400
transform 1 0 45024 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1963
timestamp 1669390400
transform 1 0 52976 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1964
timestamp 1669390400
transform 1 0 60928 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1965
timestamp 1669390400
transform 1 0 68880 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1966
timestamp 1669390400
transform 1 0 76832 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1967
timestamp 1669390400
transform 1 0 84784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1968
timestamp 1669390400
transform 1 0 92736 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1969
timestamp 1669390400
transform 1 0 100688 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1970
timestamp 1669390400
transform 1 0 108640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1971
timestamp 1669390400
transform 1 0 116592 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1972
timestamp 1669390400
transform 1 0 9296 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1973
timestamp 1669390400
transform 1 0 17248 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1974
timestamp 1669390400
transform 1 0 25200 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1975
timestamp 1669390400
transform 1 0 33152 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1976
timestamp 1669390400
transform 1 0 41104 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1977
timestamp 1669390400
transform 1 0 49056 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1978
timestamp 1669390400
transform 1 0 57008 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1979
timestamp 1669390400
transform 1 0 64960 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1980
timestamp 1669390400
transform 1 0 72912 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1981
timestamp 1669390400
transform 1 0 80864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1982
timestamp 1669390400
transform 1 0 88816 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1983
timestamp 1669390400
transform 1 0 96768 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1984
timestamp 1669390400
transform 1 0 104720 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1985
timestamp 1669390400
transform 1 0 112672 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1986
timestamp 1669390400
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1987
timestamp 1669390400
transform 1 0 13216 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1988
timestamp 1669390400
transform 1 0 21168 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1989
timestamp 1669390400
transform 1 0 29120 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1990
timestamp 1669390400
transform 1 0 37072 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1991
timestamp 1669390400
transform 1 0 45024 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1992
timestamp 1669390400
transform 1 0 52976 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1993
timestamp 1669390400
transform 1 0 60928 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1994
timestamp 1669390400
transform 1 0 68880 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1995
timestamp 1669390400
transform 1 0 76832 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1996
timestamp 1669390400
transform 1 0 84784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1997
timestamp 1669390400
transform 1 0 92736 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1998
timestamp 1669390400
transform 1 0 100688 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1999
timestamp 1669390400
transform 1 0 108640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2000
timestamp 1669390400
transform 1 0 116592 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2001
timestamp 1669390400
transform 1 0 9296 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2002
timestamp 1669390400
transform 1 0 17248 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2003
timestamp 1669390400
transform 1 0 25200 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2004
timestamp 1669390400
transform 1 0 33152 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2005
timestamp 1669390400
transform 1 0 41104 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2006
timestamp 1669390400
transform 1 0 49056 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2007
timestamp 1669390400
transform 1 0 57008 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2008
timestamp 1669390400
transform 1 0 64960 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2009
timestamp 1669390400
transform 1 0 72912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2010
timestamp 1669390400
transform 1 0 80864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2011
timestamp 1669390400
transform 1 0 88816 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2012
timestamp 1669390400
transform 1 0 96768 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2013
timestamp 1669390400
transform 1 0 104720 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2014
timestamp 1669390400
transform 1 0 112672 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2015
timestamp 1669390400
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2016
timestamp 1669390400
transform 1 0 13216 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2017
timestamp 1669390400
transform 1 0 21168 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2018
timestamp 1669390400
transform 1 0 29120 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2019
timestamp 1669390400
transform 1 0 37072 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2020
timestamp 1669390400
transform 1 0 45024 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2021
timestamp 1669390400
transform 1 0 52976 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2022
timestamp 1669390400
transform 1 0 60928 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2023
timestamp 1669390400
transform 1 0 68880 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2024
timestamp 1669390400
transform 1 0 76832 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2025
timestamp 1669390400
transform 1 0 84784 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2026
timestamp 1669390400
transform 1 0 92736 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2027
timestamp 1669390400
transform 1 0 100688 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2028
timestamp 1669390400
transform 1 0 108640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2029
timestamp 1669390400
transform 1 0 116592 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2030
timestamp 1669390400
transform 1 0 9296 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2031
timestamp 1669390400
transform 1 0 17248 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2032
timestamp 1669390400
transform 1 0 25200 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2033
timestamp 1669390400
transform 1 0 33152 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2034
timestamp 1669390400
transform 1 0 41104 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2035
timestamp 1669390400
transform 1 0 49056 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2036
timestamp 1669390400
transform 1 0 57008 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2037
timestamp 1669390400
transform 1 0 64960 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2038
timestamp 1669390400
transform 1 0 72912 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2039
timestamp 1669390400
transform 1 0 80864 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2040
timestamp 1669390400
transform 1 0 88816 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2041
timestamp 1669390400
transform 1 0 96768 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2042
timestamp 1669390400
transform 1 0 104720 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2043
timestamp 1669390400
transform 1 0 112672 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2044
timestamp 1669390400
transform 1 0 5264 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2045
timestamp 1669390400
transform 1 0 13216 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2046
timestamp 1669390400
transform 1 0 21168 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2047
timestamp 1669390400
transform 1 0 29120 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2048
timestamp 1669390400
transform 1 0 37072 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2049
timestamp 1669390400
transform 1 0 45024 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2050
timestamp 1669390400
transform 1 0 52976 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2051
timestamp 1669390400
transform 1 0 60928 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2052
timestamp 1669390400
transform 1 0 68880 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2053
timestamp 1669390400
transform 1 0 76832 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2054
timestamp 1669390400
transform 1 0 84784 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2055
timestamp 1669390400
transform 1 0 92736 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2056
timestamp 1669390400
transform 1 0 100688 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2057
timestamp 1669390400
transform 1 0 108640 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2058
timestamp 1669390400
transform 1 0 116592 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2059
timestamp 1669390400
transform 1 0 9296 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2060
timestamp 1669390400
transform 1 0 17248 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2061
timestamp 1669390400
transform 1 0 25200 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2062
timestamp 1669390400
transform 1 0 33152 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2063
timestamp 1669390400
transform 1 0 41104 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2064
timestamp 1669390400
transform 1 0 49056 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2065
timestamp 1669390400
transform 1 0 57008 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2066
timestamp 1669390400
transform 1 0 64960 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2067
timestamp 1669390400
transform 1 0 72912 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2068
timestamp 1669390400
transform 1 0 80864 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2069
timestamp 1669390400
transform 1 0 88816 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2070
timestamp 1669390400
transform 1 0 96768 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2071
timestamp 1669390400
transform 1 0 104720 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2072
timestamp 1669390400
transform 1 0 112672 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2073
timestamp 1669390400
transform 1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2074
timestamp 1669390400
transform 1 0 13216 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2075
timestamp 1669390400
transform 1 0 21168 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2076
timestamp 1669390400
transform 1 0 29120 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2077
timestamp 1669390400
transform 1 0 37072 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2078
timestamp 1669390400
transform 1 0 45024 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2079
timestamp 1669390400
transform 1 0 52976 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2080
timestamp 1669390400
transform 1 0 60928 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2081
timestamp 1669390400
transform 1 0 68880 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2082
timestamp 1669390400
transform 1 0 76832 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2083
timestamp 1669390400
transform 1 0 84784 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2084
timestamp 1669390400
transform 1 0 92736 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2085
timestamp 1669390400
transform 1 0 100688 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2086
timestamp 1669390400
transform 1 0 108640 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2087
timestamp 1669390400
transform 1 0 116592 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2088
timestamp 1669390400
transform 1 0 9296 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2089
timestamp 1669390400
transform 1 0 17248 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2090
timestamp 1669390400
transform 1 0 25200 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2091
timestamp 1669390400
transform 1 0 33152 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2092
timestamp 1669390400
transform 1 0 41104 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2093
timestamp 1669390400
transform 1 0 49056 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2094
timestamp 1669390400
transform 1 0 57008 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2095
timestamp 1669390400
transform 1 0 64960 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2096
timestamp 1669390400
transform 1 0 72912 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2097
timestamp 1669390400
transform 1 0 80864 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2098
timestamp 1669390400
transform 1 0 88816 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2099
timestamp 1669390400
transform 1 0 96768 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2100
timestamp 1669390400
transform 1 0 104720 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2101
timestamp 1669390400
transform 1 0 112672 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2102
timestamp 1669390400
transform 1 0 5264 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2103
timestamp 1669390400
transform 1 0 13216 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2104
timestamp 1669390400
transform 1 0 21168 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2105
timestamp 1669390400
transform 1 0 29120 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2106
timestamp 1669390400
transform 1 0 37072 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2107
timestamp 1669390400
transform 1 0 45024 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2108
timestamp 1669390400
transform 1 0 52976 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2109
timestamp 1669390400
transform 1 0 60928 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2110
timestamp 1669390400
transform 1 0 68880 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2111
timestamp 1669390400
transform 1 0 76832 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2112
timestamp 1669390400
transform 1 0 84784 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2113
timestamp 1669390400
transform 1 0 92736 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2114
timestamp 1669390400
transform 1 0 100688 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2115
timestamp 1669390400
transform 1 0 108640 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2116
timestamp 1669390400
transform 1 0 116592 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2117
timestamp 1669390400
transform 1 0 9296 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2118
timestamp 1669390400
transform 1 0 17248 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2119
timestamp 1669390400
transform 1 0 25200 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2120
timestamp 1669390400
transform 1 0 33152 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2121
timestamp 1669390400
transform 1 0 41104 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2122
timestamp 1669390400
transform 1 0 49056 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2123
timestamp 1669390400
transform 1 0 57008 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2124
timestamp 1669390400
transform 1 0 64960 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2125
timestamp 1669390400
transform 1 0 72912 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2126
timestamp 1669390400
transform 1 0 80864 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2127
timestamp 1669390400
transform 1 0 88816 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2128
timestamp 1669390400
transform 1 0 96768 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2129
timestamp 1669390400
transform 1 0 104720 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2130
timestamp 1669390400
transform 1 0 112672 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2131
timestamp 1669390400
transform 1 0 5264 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2132
timestamp 1669390400
transform 1 0 13216 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2133
timestamp 1669390400
transform 1 0 21168 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2134
timestamp 1669390400
transform 1 0 29120 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2135
timestamp 1669390400
transform 1 0 37072 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2136
timestamp 1669390400
transform 1 0 45024 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2137
timestamp 1669390400
transform 1 0 52976 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2138
timestamp 1669390400
transform 1 0 60928 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2139
timestamp 1669390400
transform 1 0 68880 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2140
timestamp 1669390400
transform 1 0 76832 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2141
timestamp 1669390400
transform 1 0 84784 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2142
timestamp 1669390400
transform 1 0 92736 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2143
timestamp 1669390400
transform 1 0 100688 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2144
timestamp 1669390400
transform 1 0 108640 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2145
timestamp 1669390400
transform 1 0 116592 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2146
timestamp 1669390400
transform 1 0 9296 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2147
timestamp 1669390400
transform 1 0 17248 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2148
timestamp 1669390400
transform 1 0 25200 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2149
timestamp 1669390400
transform 1 0 33152 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2150
timestamp 1669390400
transform 1 0 41104 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2151
timestamp 1669390400
transform 1 0 49056 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2152
timestamp 1669390400
transform 1 0 57008 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2153
timestamp 1669390400
transform 1 0 64960 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2154
timestamp 1669390400
transform 1 0 72912 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2155
timestamp 1669390400
transform 1 0 80864 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2156
timestamp 1669390400
transform 1 0 88816 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2157
timestamp 1669390400
transform 1 0 96768 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2158
timestamp 1669390400
transform 1 0 104720 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2159
timestamp 1669390400
transform 1 0 112672 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2160
timestamp 1669390400
transform 1 0 5264 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2161
timestamp 1669390400
transform 1 0 13216 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2162
timestamp 1669390400
transform 1 0 21168 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2163
timestamp 1669390400
transform 1 0 29120 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2164
timestamp 1669390400
transform 1 0 37072 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2165
timestamp 1669390400
transform 1 0 45024 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2166
timestamp 1669390400
transform 1 0 52976 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2167
timestamp 1669390400
transform 1 0 60928 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2168
timestamp 1669390400
transform 1 0 68880 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2169
timestamp 1669390400
transform 1 0 76832 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2170
timestamp 1669390400
transform 1 0 84784 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2171
timestamp 1669390400
transform 1 0 92736 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2172
timestamp 1669390400
transform 1 0 100688 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2173
timestamp 1669390400
transform 1 0 108640 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2174
timestamp 1669390400
transform 1 0 116592 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2175
timestamp 1669390400
transform 1 0 9296 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2176
timestamp 1669390400
transform 1 0 17248 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2177
timestamp 1669390400
transform 1 0 25200 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2178
timestamp 1669390400
transform 1 0 33152 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2179
timestamp 1669390400
transform 1 0 41104 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2180
timestamp 1669390400
transform 1 0 49056 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2181
timestamp 1669390400
transform 1 0 57008 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2182
timestamp 1669390400
transform 1 0 64960 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2183
timestamp 1669390400
transform 1 0 72912 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2184
timestamp 1669390400
transform 1 0 80864 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2185
timestamp 1669390400
transform 1 0 88816 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2186
timestamp 1669390400
transform 1 0 96768 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2187
timestamp 1669390400
transform 1 0 104720 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2188
timestamp 1669390400
transform 1 0 112672 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2189
timestamp 1669390400
transform 1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2190
timestamp 1669390400
transform 1 0 13216 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2191
timestamp 1669390400
transform 1 0 21168 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2192
timestamp 1669390400
transform 1 0 29120 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2193
timestamp 1669390400
transform 1 0 37072 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2194
timestamp 1669390400
transform 1 0 45024 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2195
timestamp 1669390400
transform 1 0 52976 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2196
timestamp 1669390400
transform 1 0 60928 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2197
timestamp 1669390400
transform 1 0 68880 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2198
timestamp 1669390400
transform 1 0 76832 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2199
timestamp 1669390400
transform 1 0 84784 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2200
timestamp 1669390400
transform 1 0 92736 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2201
timestamp 1669390400
transform 1 0 100688 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2202
timestamp 1669390400
transform 1 0 108640 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2203
timestamp 1669390400
transform 1 0 116592 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2204
timestamp 1669390400
transform 1 0 9296 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2205
timestamp 1669390400
transform 1 0 17248 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2206
timestamp 1669390400
transform 1 0 25200 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2207
timestamp 1669390400
transform 1 0 33152 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2208
timestamp 1669390400
transform 1 0 41104 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2209
timestamp 1669390400
transform 1 0 49056 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2210
timestamp 1669390400
transform 1 0 57008 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2211
timestamp 1669390400
transform 1 0 64960 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2212
timestamp 1669390400
transform 1 0 72912 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2213
timestamp 1669390400
transform 1 0 80864 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2214
timestamp 1669390400
transform 1 0 88816 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2215
timestamp 1669390400
transform 1 0 96768 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2216
timestamp 1669390400
transform 1 0 104720 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2217
timestamp 1669390400
transform 1 0 112672 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2218
timestamp 1669390400
transform 1 0 5264 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2219
timestamp 1669390400
transform 1 0 13216 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2220
timestamp 1669390400
transform 1 0 21168 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2221
timestamp 1669390400
transform 1 0 29120 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2222
timestamp 1669390400
transform 1 0 37072 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2223
timestamp 1669390400
transform 1 0 45024 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2224
timestamp 1669390400
transform 1 0 52976 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2225
timestamp 1669390400
transform 1 0 60928 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2226
timestamp 1669390400
transform 1 0 68880 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2227
timestamp 1669390400
transform 1 0 76832 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2228
timestamp 1669390400
transform 1 0 84784 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2229
timestamp 1669390400
transform 1 0 92736 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2230
timestamp 1669390400
transform 1 0 100688 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2231
timestamp 1669390400
transform 1 0 108640 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2232
timestamp 1669390400
transform 1 0 116592 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2233
timestamp 1669390400
transform 1 0 9296 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2234
timestamp 1669390400
transform 1 0 17248 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2235
timestamp 1669390400
transform 1 0 25200 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2236
timestamp 1669390400
transform 1 0 33152 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2237
timestamp 1669390400
transform 1 0 41104 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2238
timestamp 1669390400
transform 1 0 49056 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2239
timestamp 1669390400
transform 1 0 57008 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2240
timestamp 1669390400
transform 1 0 64960 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2241
timestamp 1669390400
transform 1 0 72912 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2242
timestamp 1669390400
transform 1 0 80864 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2243
timestamp 1669390400
transform 1 0 88816 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2244
timestamp 1669390400
transform 1 0 96768 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2245
timestamp 1669390400
transform 1 0 104720 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2246
timestamp 1669390400
transform 1 0 112672 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2247
timestamp 1669390400
transform 1 0 5264 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2248
timestamp 1669390400
transform 1 0 13216 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2249
timestamp 1669390400
transform 1 0 21168 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2250
timestamp 1669390400
transform 1 0 29120 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2251
timestamp 1669390400
transform 1 0 37072 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2252
timestamp 1669390400
transform 1 0 45024 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2253
timestamp 1669390400
transform 1 0 52976 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2254
timestamp 1669390400
transform 1 0 60928 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2255
timestamp 1669390400
transform 1 0 68880 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2256
timestamp 1669390400
transform 1 0 76832 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2257
timestamp 1669390400
transform 1 0 84784 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2258
timestamp 1669390400
transform 1 0 92736 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2259
timestamp 1669390400
transform 1 0 100688 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2260
timestamp 1669390400
transform 1 0 108640 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2261
timestamp 1669390400
transform 1 0 116592 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2262
timestamp 1669390400
transform 1 0 9296 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2263
timestamp 1669390400
transform 1 0 17248 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2264
timestamp 1669390400
transform 1 0 25200 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2265
timestamp 1669390400
transform 1 0 33152 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2266
timestamp 1669390400
transform 1 0 41104 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2267
timestamp 1669390400
transform 1 0 49056 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2268
timestamp 1669390400
transform 1 0 57008 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2269
timestamp 1669390400
transform 1 0 64960 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2270
timestamp 1669390400
transform 1 0 72912 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2271
timestamp 1669390400
transform 1 0 80864 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2272
timestamp 1669390400
transform 1 0 88816 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2273
timestamp 1669390400
transform 1 0 96768 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2274
timestamp 1669390400
transform 1 0 104720 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2275
timestamp 1669390400
transform 1 0 112672 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2276
timestamp 1669390400
transform 1 0 5264 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2277
timestamp 1669390400
transform 1 0 13216 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2278
timestamp 1669390400
transform 1 0 21168 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2279
timestamp 1669390400
transform 1 0 29120 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2280
timestamp 1669390400
transform 1 0 37072 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2281
timestamp 1669390400
transform 1 0 45024 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2282
timestamp 1669390400
transform 1 0 52976 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2283
timestamp 1669390400
transform 1 0 60928 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2284
timestamp 1669390400
transform 1 0 68880 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2285
timestamp 1669390400
transform 1 0 76832 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2286
timestamp 1669390400
transform 1 0 84784 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2287
timestamp 1669390400
transform 1 0 92736 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2288
timestamp 1669390400
transform 1 0 100688 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2289
timestamp 1669390400
transform 1 0 108640 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2290
timestamp 1669390400
transform 1 0 116592 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2291
timestamp 1669390400
transform 1 0 9296 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2292
timestamp 1669390400
transform 1 0 17248 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2293
timestamp 1669390400
transform 1 0 25200 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2294
timestamp 1669390400
transform 1 0 33152 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2295
timestamp 1669390400
transform 1 0 41104 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2296
timestamp 1669390400
transform 1 0 49056 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2297
timestamp 1669390400
transform 1 0 57008 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2298
timestamp 1669390400
transform 1 0 64960 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2299
timestamp 1669390400
transform 1 0 72912 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2300
timestamp 1669390400
transform 1 0 80864 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2301
timestamp 1669390400
transform 1 0 88816 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2302
timestamp 1669390400
transform 1 0 96768 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2303
timestamp 1669390400
transform 1 0 104720 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2304
timestamp 1669390400
transform 1 0 112672 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2305
timestamp 1669390400
transform 1 0 5264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2306
timestamp 1669390400
transform 1 0 13216 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2307
timestamp 1669390400
transform 1 0 21168 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2308
timestamp 1669390400
transform 1 0 29120 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2309
timestamp 1669390400
transform 1 0 37072 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2310
timestamp 1669390400
transform 1 0 45024 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2311
timestamp 1669390400
transform 1 0 52976 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2312
timestamp 1669390400
transform 1 0 60928 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2313
timestamp 1669390400
transform 1 0 68880 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2314
timestamp 1669390400
transform 1 0 76832 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2315
timestamp 1669390400
transform 1 0 84784 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2316
timestamp 1669390400
transform 1 0 92736 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2317
timestamp 1669390400
transform 1 0 100688 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2318
timestamp 1669390400
transform 1 0 108640 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2319
timestamp 1669390400
transform 1 0 116592 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2320
timestamp 1669390400
transform 1 0 9296 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2321
timestamp 1669390400
transform 1 0 17248 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2322
timestamp 1669390400
transform 1 0 25200 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2323
timestamp 1669390400
transform 1 0 33152 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2324
timestamp 1669390400
transform 1 0 41104 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2325
timestamp 1669390400
transform 1 0 49056 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2326
timestamp 1669390400
transform 1 0 57008 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2327
timestamp 1669390400
transform 1 0 64960 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2328
timestamp 1669390400
transform 1 0 72912 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2329
timestamp 1669390400
transform 1 0 80864 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2330
timestamp 1669390400
transform 1 0 88816 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2331
timestamp 1669390400
transform 1 0 96768 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2332
timestamp 1669390400
transform 1 0 104720 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2333
timestamp 1669390400
transform 1 0 112672 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2334
timestamp 1669390400
transform 1 0 5264 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2335
timestamp 1669390400
transform 1 0 13216 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2336
timestamp 1669390400
transform 1 0 21168 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2337
timestamp 1669390400
transform 1 0 29120 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2338
timestamp 1669390400
transform 1 0 37072 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2339
timestamp 1669390400
transform 1 0 45024 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2340
timestamp 1669390400
transform 1 0 52976 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2341
timestamp 1669390400
transform 1 0 60928 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2342
timestamp 1669390400
transform 1 0 68880 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2343
timestamp 1669390400
transform 1 0 76832 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2344
timestamp 1669390400
transform 1 0 84784 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2345
timestamp 1669390400
transform 1 0 92736 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2346
timestamp 1669390400
transform 1 0 100688 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2347
timestamp 1669390400
transform 1 0 108640 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2348
timestamp 1669390400
transform 1 0 116592 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2349
timestamp 1669390400
transform 1 0 9296 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2350
timestamp 1669390400
transform 1 0 17248 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2351
timestamp 1669390400
transform 1 0 25200 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2352
timestamp 1669390400
transform 1 0 33152 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2353
timestamp 1669390400
transform 1 0 41104 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2354
timestamp 1669390400
transform 1 0 49056 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2355
timestamp 1669390400
transform 1 0 57008 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2356
timestamp 1669390400
transform 1 0 64960 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2357
timestamp 1669390400
transform 1 0 72912 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2358
timestamp 1669390400
transform 1 0 80864 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2359
timestamp 1669390400
transform 1 0 88816 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2360
timestamp 1669390400
transform 1 0 96768 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2361
timestamp 1669390400
transform 1 0 104720 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2362
timestamp 1669390400
transform 1 0 112672 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2363
timestamp 1669390400
transform 1 0 5264 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2364
timestamp 1669390400
transform 1 0 13216 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2365
timestamp 1669390400
transform 1 0 21168 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2366
timestamp 1669390400
transform 1 0 29120 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2367
timestamp 1669390400
transform 1 0 37072 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2368
timestamp 1669390400
transform 1 0 45024 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2369
timestamp 1669390400
transform 1 0 52976 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2370
timestamp 1669390400
transform 1 0 60928 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2371
timestamp 1669390400
transform 1 0 68880 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2372
timestamp 1669390400
transform 1 0 76832 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2373
timestamp 1669390400
transform 1 0 84784 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2374
timestamp 1669390400
transform 1 0 92736 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2375
timestamp 1669390400
transform 1 0 100688 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2376
timestamp 1669390400
transform 1 0 108640 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2377
timestamp 1669390400
transform 1 0 116592 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2378
timestamp 1669390400
transform 1 0 9296 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2379
timestamp 1669390400
transform 1 0 17248 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2380
timestamp 1669390400
transform 1 0 25200 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2381
timestamp 1669390400
transform 1 0 33152 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2382
timestamp 1669390400
transform 1 0 41104 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2383
timestamp 1669390400
transform 1 0 49056 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2384
timestamp 1669390400
transform 1 0 57008 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2385
timestamp 1669390400
transform 1 0 64960 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2386
timestamp 1669390400
transform 1 0 72912 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2387
timestamp 1669390400
transform 1 0 80864 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2388
timestamp 1669390400
transform 1 0 88816 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2389
timestamp 1669390400
transform 1 0 96768 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2390
timestamp 1669390400
transform 1 0 104720 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2391
timestamp 1669390400
transform 1 0 112672 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2392
timestamp 1669390400
transform 1 0 5264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2393
timestamp 1669390400
transform 1 0 9184 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2394
timestamp 1669390400
transform 1 0 13104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2395
timestamp 1669390400
transform 1 0 17024 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2396
timestamp 1669390400
transform 1 0 20944 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2397
timestamp 1669390400
transform 1 0 24864 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2398
timestamp 1669390400
transform 1 0 28784 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2399
timestamp 1669390400
transform 1 0 32704 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2400
timestamp 1669390400
transform 1 0 36624 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2401
timestamp 1669390400
transform 1 0 40544 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2402
timestamp 1669390400
transform 1 0 44464 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2403
timestamp 1669390400
transform 1 0 48384 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2404
timestamp 1669390400
transform 1 0 52304 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2405
timestamp 1669390400
transform 1 0 56224 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2406
timestamp 1669390400
transform 1 0 60144 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2407
timestamp 1669390400
transform 1 0 64064 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2408
timestamp 1669390400
transform 1 0 67984 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2409
timestamp 1669390400
transform 1 0 71904 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2410
timestamp 1669390400
transform 1 0 75824 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2411
timestamp 1669390400
transform 1 0 79744 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2412
timestamp 1669390400
transform 1 0 83664 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2413
timestamp 1669390400
transform 1 0 87584 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2414
timestamp 1669390400
transform 1 0 91504 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2415
timestamp 1669390400
transform 1 0 95424 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2416
timestamp 1669390400
transform 1 0 99344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2417
timestamp 1669390400
transform 1 0 103264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2418
timestamp 1669390400
transform 1 0 107184 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2419
timestamp 1669390400
transform 1 0 111104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2420
timestamp 1669390400
transform 1 0 115024 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _298_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 63952 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _299_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 62496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _300_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38192 0 1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _301_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41552 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1669390400
transform 1 0 52752 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _303_
timestamp 1669390400
transform 1 0 53312 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _304_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 63056 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _305_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 60144 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _306_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 61264 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _307_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 47376 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _308_
timestamp 1669390400
transform 1 0 70784 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _309_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 48160 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _310_
timestamp 1669390400
transform 1 0 47376 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _311_
timestamp 1669390400
transform -1 0 47936 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _312_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 46704 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _313_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 90944 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _314_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 91616 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _315_
timestamp 1669390400
transform 1 0 115808 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _316_
timestamp 1669390400
transform -1 0 116480 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _317_
timestamp 1669390400
transform 1 0 45808 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _318_
timestamp 1669390400
transform 1 0 44016 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _319_
timestamp 1669390400
transform 1 0 45808 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _320_
timestamp 1669390400
transform 1 0 45360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _321_
timestamp 1669390400
transform 1 0 47376 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _322_
timestamp 1669390400
transform 1 0 45472 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_
timestamp 1669390400
transform 1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _324_
timestamp 1669390400
transform 1 0 114800 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1669390400
transform 1 0 113904 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _326_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 69216 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _327_
timestamp 1669390400
transform 1 0 71904 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _328_
timestamp 1669390400
transform 1 0 69664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _329_
timestamp 1669390400
transform 1 0 77616 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1669390400
transform 1 0 77280 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _331_
timestamp 1669390400
transform 1 0 74592 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _332_
timestamp 1669390400
transform 1 0 74592 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _333_
timestamp 1669390400
transform 1 0 65184 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _334_
timestamp 1669390400
transform 1 0 67200 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _335_
timestamp 1669390400
transform 1 0 65968 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _336_
timestamp 1669390400
transform 1 0 45472 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1669390400
transform 1 0 45360 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _338_
timestamp 1669390400
transform -1 0 117824 0 -1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _339_
timestamp 1669390400
transform -1 0 117600 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _340_
timestamp 1669390400
transform 1 0 71120 0 -1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _341_
timestamp 1669390400
transform 1 0 71568 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _342_
timestamp 1669390400
transform 1 0 53536 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _343_
timestamp 1669390400
transform 1 0 71904 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _344_
timestamp 1669390400
transform 1 0 70784 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _345_
timestamp 1669390400
transform -1 0 68208 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _346_
timestamp 1669390400
transform 1 0 70336 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _347_
timestamp 1669390400
transform 1 0 69216 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _348_
timestamp 1669390400
transform 1 0 45808 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1669390400
transform 1 0 45584 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _350_
timestamp 1669390400
transform 1 0 53984 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _351_
timestamp 1669390400
transform 1 0 53312 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _352_
timestamp 1669390400
transform 1 0 78288 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1669390400
transform 1 0 77392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _354_
timestamp 1669390400
transform 1 0 45472 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1669390400
transform 1 0 45360 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _356_
timestamp 1669390400
transform 1 0 46144 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _357_
timestamp 1669390400
transform 1 0 45696 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _358_
timestamp 1669390400
transform 1 0 45360 0 1 64288
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1669390400
transform 1 0 45360 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _360_
timestamp 1669390400
transform -1 0 49168 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _361_
timestamp 1669390400
transform -1 0 50064 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _362_
timestamp 1669390400
transform 1 0 47712 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _363_
timestamp 1669390400
transform -1 0 52304 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _364_
timestamp 1669390400
transform -1 0 48384 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _365_
timestamp 1669390400
transform 1 0 46592 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _366_
timestamp 1669390400
transform 1 0 47824 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _367_
timestamp 1669390400
transform 1 0 47264 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _368_
timestamp 1669390400
transform -1 0 50176 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _369_
timestamp 1669390400
transform -1 0 48048 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _370_
timestamp 1669390400
transform 1 0 47152 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _371_
timestamp 1669390400
transform 1 0 61264 0 1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1669390400
transform 1 0 61264 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _373_
timestamp 1669390400
transform 1 0 49392 0 -1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1669390400
transform 1 0 48160 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _375_
timestamp 1669390400
transform 1 0 61488 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _376_
timestamp 1669390400
transform 1 0 61376 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _377_
timestamp 1669390400
transform -1 0 71232 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _378_
timestamp 1669390400
transform 1 0 73248 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _379_
timestamp 1669390400
transform 1 0 71568 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _380_
timestamp 1669390400
transform -1 0 68880 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _381_
timestamp 1669390400
transform 1 0 50288 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _382_
timestamp 1669390400
transform 1 0 49952 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _383_
timestamp 1669390400
transform 1 0 70672 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _384_
timestamp 1669390400
transform 1 0 73248 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _385_
timestamp 1669390400
transform 1 0 71680 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _386_
timestamp 1669390400
transform -1 0 56672 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _387_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54096 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _388_
timestamp 1669390400
transform 1 0 67424 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _389_
timestamp 1669390400
transform 1 0 62832 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _390_
timestamp 1669390400
transform 1 0 65632 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _391_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 66640 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _392_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 62608 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _393_
timestamp 1669390400
transform -1 0 60144 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _394_
timestamp 1669390400
transform -1 0 55104 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _395_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55328 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _396_
timestamp 1669390400
transform -1 0 54208 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _397_
timestamp 1669390400
transform -1 0 56560 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _398_
timestamp 1669390400
transform -1 0 54432 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _399_
timestamp 1669390400
transform 1 0 41440 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _400_
timestamp 1669390400
transform -1 0 41104 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _401_
timestamp 1669390400
transform 1 0 67872 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _402_
timestamp 1669390400
transform -1 0 52864 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _403_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _404_
timestamp 1669390400
transform 1 0 54208 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _405_
timestamp 1669390400
transform 1 0 60704 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _406_
timestamp 1669390400
transform 1 0 62048 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _407_
timestamp 1669390400
transform -1 0 58800 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _408_
timestamp 1669390400
transform -1 0 54544 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _409_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 59136 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _410_
timestamp 1669390400
transform 1 0 61264 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _411_
timestamp 1669390400
transform 1 0 67648 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _412_
timestamp 1669390400
transform 1 0 61040 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _413_
timestamp 1669390400
transform -1 0 58464 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _414_
timestamp 1669390400
transform 1 0 59696 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _415_
timestamp 1669390400
transform 1 0 58912 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _416_
timestamp 1669390400
transform -1 0 43568 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _417_
timestamp 1669390400
transform 1 0 63392 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _418_
timestamp 1669390400
transform -1 0 58464 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _419_
timestamp 1669390400
transform -1 0 59808 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _420_
timestamp 1669390400
transform -1 0 60368 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _421_
timestamp 1669390400
transform 1 0 59696 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _422_
timestamp 1669390400
transform -1 0 58576 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _423_
timestamp 1669390400
transform -1 0 59248 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _424_
timestamp 1669390400
transform 1 0 58800 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _425_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 58912 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _426_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56896 0 -1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _427_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 59024 0 1 50176
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _428_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 59584 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _429_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 64848 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _430_
timestamp 1669390400
transform 1 0 61264 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _431_
timestamp 1669390400
transform 1 0 63840 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _432_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54544 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _433_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54880 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _434_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55440 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _435_
timestamp 1669390400
transform -1 0 56224 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _436_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 64512 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _437_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 62272 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _438_
timestamp 1669390400
transform -1 0 63504 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _439_
timestamp 1669390400
transform 1 0 64176 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _440_
timestamp 1669390400
transform 1 0 63840 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _441_
timestamp 1669390400
transform 1 0 61152 0 -1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _442_
timestamp 1669390400
transform -1 0 60928 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _443_
timestamp 1669390400
transform -1 0 59248 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _444_
timestamp 1669390400
transform -1 0 59248 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _445_
timestamp 1669390400
transform 1 0 59472 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _446_
timestamp 1669390400
transform -1 0 58912 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _447_
timestamp 1669390400
transform -1 0 58016 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _448_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 62832 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _449_
timestamp 1669390400
transform -1 0 59248 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _450_
timestamp 1669390400
transform 1 0 57344 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _451_
timestamp 1669390400
transform 1 0 57568 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _452_
timestamp 1669390400
transform 1 0 58128 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _453_
timestamp 1669390400
transform -1 0 59808 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _454_
timestamp 1669390400
transform 1 0 58688 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _455_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 60368 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _456_
timestamp 1669390400
transform 1 0 61264 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _457_
timestamp 1669390400
transform 1 0 58464 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _458_
timestamp 1669390400
transform 1 0 61264 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _459_
timestamp 1669390400
transform -1 0 63840 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _460_
timestamp 1669390400
transform 1 0 62496 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _461_
timestamp 1669390400
transform 1 0 63728 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _462_
timestamp 1669390400
transform -1 0 64176 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _463_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 62272 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _464_
timestamp 1669390400
transform 1 0 63280 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _465_
timestamp 1669390400
transform -1 0 64848 0 -1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _466_
timestamp 1669390400
transform 1 0 65184 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _467_
timestamp 1669390400
transform -1 0 64064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _468_
timestamp 1669390400
transform 1 0 54320 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _469_
timestamp 1669390400
transform 1 0 57344 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _470_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 57232 0 1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _471_
timestamp 1669390400
transform -1 0 65968 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _472_
timestamp 1669390400
transform -1 0 64176 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _473_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56560 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _474_
timestamp 1669390400
transform 1 0 62496 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _475_
timestamp 1669390400
transform 1 0 65296 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _476_
timestamp 1669390400
transform 1 0 63504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _477_
timestamp 1669390400
transform -1 0 65856 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _478_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 64400 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _479_
timestamp 1669390400
transform -1 0 63392 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _480_
timestamp 1669390400
transform -1 0 62384 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _481_
timestamp 1669390400
transform -1 0 60032 0 -1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _482_
timestamp 1669390400
transform 1 0 61264 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _483_
timestamp 1669390400
transform -1 0 64624 0 1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _484_
timestamp 1669390400
transform 1 0 62048 0 -1 65856
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _485_
timestamp 1669390400
transform 1 0 63168 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _486_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 63616 0 1 62720
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _487_
timestamp 1669390400
transform -1 0 56112 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _488_
timestamp 1669390400
transform 1 0 54320 0 -1 62720
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _489_
timestamp 1669390400
transform -1 0 54544 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _490_
timestamp 1669390400
transform -1 0 56336 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _491_
timestamp 1669390400
transform 1 0 54544 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _492_
timestamp 1669390400
transform 1 0 54432 0 1 65856
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _493_
timestamp 1669390400
transform -1 0 54208 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _494_
timestamp 1669390400
transform 1 0 56112 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _495_
timestamp 1669390400
transform 1 0 56112 0 1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _496_
timestamp 1669390400
transform 1 0 56224 0 1 65856
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _497_
timestamp 1669390400
transform 1 0 58016 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _498_
timestamp 1669390400
transform -1 0 59696 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _499_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54320 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _500_
timestamp 1669390400
transform 1 0 55440 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _501_
timestamp 1669390400
transform 1 0 53648 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _502_
timestamp 1669390400
transform 1 0 54768 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _503_
timestamp 1669390400
transform -1 0 56000 0 1 59584
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _504_
timestamp 1669390400
transform -1 0 54544 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _505_
timestamp 1669390400
transform 1 0 57344 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _506_
timestamp 1669390400
transform -1 0 59360 0 1 62720
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _507_
timestamp 1669390400
transform 1 0 58016 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _508_
timestamp 1669390400
transform -1 0 59808 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1669390400
transform -1 0 61824 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _510_
timestamp 1669390400
transform -1 0 59136 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _511_
timestamp 1669390400
transform 1 0 57344 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _512_
timestamp 1669390400
transform 1 0 56672 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _513_
timestamp 1669390400
transform 1 0 57344 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _514_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 58464 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _515_
timestamp 1669390400
transform -1 0 58912 0 -1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _516_
timestamp 1669390400
transform 1 0 59136 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _517_
timestamp 1669390400
transform 1 0 52752 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _518_
timestamp 1669390400
transform -1 0 56672 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _519_
timestamp 1669390400
transform 1 0 57120 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _520_
timestamp 1669390400
transform 1 0 57344 0 -1 58016
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _521_
timestamp 1669390400
transform -1 0 54096 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _522_
timestamp 1669390400
transform -1 0 55552 0 -1 56448
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _523_
timestamp 1669390400
transform 1 0 54880 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _524_
timestamp 1669390400
transform 1 0 60592 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _525_
timestamp 1669390400
transform -1 0 63280 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _526_
timestamp 1669390400
transform 1 0 63504 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _527_
timestamp 1669390400
transform 1 0 63728 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _528_
timestamp 1669390400
transform 1 0 51408 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _529_
timestamp 1669390400
transform -1 0 51744 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _530_
timestamp 1669390400
transform 1 0 51632 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _531_
timestamp 1669390400
transform -1 0 50736 0 -1 56448
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _532_
timestamp 1669390400
transform -1 0 50176 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _533_
timestamp 1669390400
transform 1 0 51296 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _534_
timestamp 1669390400
transform 1 0 51184 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _535_
timestamp 1669390400
transform 1 0 53312 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _536_
timestamp 1669390400
transform 1 0 51744 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _537_
timestamp 1669390400
transform 1 0 51856 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _538_
timestamp 1669390400
transform 1 0 52192 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _539_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _540_
timestamp 1669390400
transform -1 0 67648 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _541_
timestamp 1669390400
transform -1 0 55552 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _542_
timestamp 1669390400
transform -1 0 51072 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _543_
timestamp 1669390400
transform 1 0 49392 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _544_
timestamp 1669390400
transform 1 0 50512 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _545_
timestamp 1669390400
transform 1 0 66528 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _546_
timestamp 1669390400
transform 1 0 50400 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _547_
timestamp 1669390400
transform 1 0 66080 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _548_
timestamp 1669390400
transform 1 0 66304 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _549_
timestamp 1669390400
transform 1 0 67760 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _550_
timestamp 1669390400
transform 1 0 54096 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _551_
timestamp 1669390400
transform -1 0 54544 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _552_
timestamp 1669390400
transform 1 0 54768 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _553_
timestamp 1669390400
transform 1 0 66416 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _554_
timestamp 1669390400
transform 1 0 66416 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _555_
timestamp 1669390400
transform -1 0 56896 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _556_
timestamp 1669390400
transform -1 0 68096 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _557_
timestamp 1669390400
transform 1 0 68320 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _558_
timestamp 1669390400
transform -1 0 51968 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _559_
timestamp 1669390400
transform -1 0 52304 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _560_
timestamp 1669390400
transform -1 0 51296 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _561_
timestamp 1669390400
transform 1 0 49392 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _562_
timestamp 1669390400
transform -1 0 54320 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _563_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 51072 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _564_
timestamp 1669390400
transform -1 0 51296 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _565_
timestamp 1669390400
transform 1 0 50960 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _566_
timestamp 1669390400
transform -1 0 50736 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _567_
timestamp 1669390400
transform -1 0 50736 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _568_
timestamp 1669390400
transform 1 0 49392 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _569_
timestamp 1669390400
transform 1 0 48048 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _570_
timestamp 1669390400
transform -1 0 50288 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _571_
timestamp 1669390400
transform 1 0 49952 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _572_
timestamp 1669390400
transform -1 0 69104 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _573_
timestamp 1669390400
transform -1 0 67648 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _574_
timestamp 1669390400
transform -1 0 50288 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _575_
timestamp 1669390400
transform -1 0 49728 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _576_
timestamp 1669390400
transform -1 0 52528 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _577_
timestamp 1669390400
transform -1 0 50848 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _578_
timestamp 1669390400
transform 1 0 49168 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _579_
timestamp 1669390400
transform 1 0 50512 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _580_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 69216 0 1 58016
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _581_
timestamp 1669390400
transform -1 0 70784 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _582_
timestamp 1669390400
transform 1 0 69216 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _583_
timestamp 1669390400
transform -1 0 70560 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _584_
timestamp 1669390400
transform 1 0 70112 0 -1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _585_
timestamp 1669390400
transform 1 0 69216 0 1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _586_
timestamp 1669390400
transform -1 0 70336 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _587_
timestamp 1669390400
transform 1 0 70672 0 1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _588_
timestamp 1669390400
transform -1 0 69104 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _589_
timestamp 1669390400
transform -1 0 69888 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _590_
timestamp 1669390400
transform -1 0 70336 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _591_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 70560 0 -1 61152
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _592_
timestamp 1669390400
transform -1 0 68768 0 1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _593_
timestamp 1669390400
transform 1 0 65744 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _594_
timestamp 1669390400
transform -1 0 68096 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _595_
timestamp 1669390400
transform 1 0 67312 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _596_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 70224 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _597_
timestamp 1669390400
transform -1 0 48608 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _598_
timestamp 1669390400
transform 1 0 91056 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _599_
timestamp 1669390400
transform 1 0 115024 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _600_
timestamp 1669390400
transform -1 0 48160 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _601_
timestamp 1669390400
transform -1 0 48608 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _602_
timestamp 1669390400
transform -1 0 47824 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _603_
timestamp 1669390400
transform 1 0 114352 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _604_
timestamp 1669390400
transform 1 0 69216 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _605_
timestamp 1669390400
transform 1 0 77504 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _606_
timestamp 1669390400
transform 1 0 74032 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _607_
timestamp 1669390400
transform 1 0 65520 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _608_
timestamp 1669390400
transform 1 0 45360 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _609_
timestamp 1669390400
transform -1 0 118272 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _610_
timestamp 1669390400
transform 1 0 71120 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _611_
timestamp 1669390400
transform 1 0 70448 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _612_
timestamp 1669390400
transform 1 0 68992 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _613_
timestamp 1669390400
transform -1 0 48160 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _614_
timestamp 1669390400
transform 1 0 53312 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _615_
timestamp 1669390400
transform 1 0 77392 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _616_
timestamp 1669390400
transform -1 0 47936 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _617_
timestamp 1669390400
transform -1 0 48048 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _618_
timestamp 1669390400
transform -1 0 47712 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _619_
timestamp 1669390400
transform -1 0 48944 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _620_
timestamp 1669390400
transform -1 0 48608 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _621_
timestamp 1669390400
transform -1 0 48944 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _622_
timestamp 1669390400
transform -1 0 48720 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _623_
timestamp 1669390400
transform 1 0 61040 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _624_
timestamp 1669390400
transform -1 0 50400 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _625_
timestamp 1669390400
transform 1 0 61264 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _626_
timestamp 1669390400
transform 1 0 71456 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _627_
timestamp 1669390400
transform -1 0 51744 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _628_
timestamp 1669390400
transform 1 0 71456 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _629_ gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 60144 0 -1 51744
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _630_
timestamp 1669390400
transform 1 0 54432 0 1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _631_
timestamp 1669390400
transform 1 0 63728 0 1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _632_
timestamp 1669390400
transform 1 0 59024 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _633_
timestamp 1669390400
transform -1 0 60480 0 1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _634_
timestamp 1669390400
transform 1 0 60816 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _635_
timestamp 1669390400
transform -1 0 67200 0 1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _636_
timestamp 1669390400
transform 1 0 65520 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _637_
timestamp 1669390400
transform -1 0 66752 0 1 59584
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _638_
timestamp 1669390400
transform -1 0 62832 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _639_
timestamp 1669390400
transform 1 0 62832 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _640_
timestamp 1669390400
transform 1 0 53312 0 1 62720
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _641_
timestamp 1669390400
transform 1 0 52416 0 -1 67424
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _642_
timestamp 1669390400
transform 1 0 57344 0 -1 67424
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _643_
timestamp 1669390400
transform -1 0 53872 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _644_
timestamp 1669390400
transform 1 0 58912 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _645_
timestamp 1669390400
transform 1 0 59808 0 -1 54880
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _646_
timestamp 1669390400
transform 1 0 53648 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _647_
timestamp 1669390400
transform 1 0 63056 0 1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _648_
timestamp 1669390400
transform 1 0 48272 0 1 56448
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _649_
timestamp 1669390400
transform 1 0 53312 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _650_
timestamp 1669390400
transform 1 0 53312 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _651_
timestamp 1669390400
transform 1 0 49616 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _652_
timestamp 1669390400
transform 1 0 67648 0 -1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _653_
timestamp 1669390400
transform 1 0 67760 0 -1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _654_
timestamp 1669390400
transform -1 0 52080 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _655_
timestamp 1669390400
transform 1 0 48160 0 1 58016
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _656_
timestamp 1669390400
transform -1 0 48944 0 -1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _657_
timestamp 1669390400
transform 1 0 50400 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _658_
timestamp 1669390400
transform 1 0 69552 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _659_
timestamp 1669390400
transform 1 0 70000 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _660_
timestamp 1669390400
transform 1 0 66528 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _703_
timestamp 1669390400
transform 1 0 3472 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _704_
timestamp 1669390400
transform -1 0 117600 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _705_
timestamp 1669390400
transform 1 0 76832 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _706_
timestamp 1669390400
transform -1 0 117600 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _707_
timestamp 1669390400
transform -1 0 4368 0 1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _708_
timestamp 1669390400
transform -1 0 117600 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _709_
timestamp 1669390400
transform 1 0 57344 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _710_
timestamp 1669390400
transform -1 0 117600 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _711_
timestamp 1669390400
transform -1 0 117600 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _712_
timestamp 1669390400
transform -1 0 117600 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _713_
timestamp 1669390400
transform -1 0 3024 0 1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _714_
timestamp 1669390400
transform -1 0 3024 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _715_
timestamp 1669390400
transform -1 0 3024 0 1 89376
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _716_
timestamp 1669390400
transform 1 0 103376 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _717_
timestamp 1669390400
transform -1 0 117600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _718_
timestamp 1669390400
transform 1 0 63392 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _719_
timestamp 1669390400
transform -1 0 3024 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _720_
timestamp 1669390400
transform 1 0 10192 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _721_
timestamp 1669390400
transform -1 0 3024 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _722_
timestamp 1669390400
transform 1 0 48272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _723_
timestamp 1669390400
transform 1 0 100688 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _724_
timestamp 1669390400
transform 1 0 10976 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _725_
timestamp 1669390400
transform -1 0 117600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _726_
timestamp 1669390400
transform 1 0 2352 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _727_
timestamp 1669390400
transform -1 0 117600 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _728_
timestamp 1669390400
transform 1 0 42224 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _729_
timestamp 1669390400
transform 1 0 99008 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _730_
timestamp 1669390400
transform -1 0 3024 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _731_
timestamp 1669390400
transform -1 0 3024 0 1 112896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _732_
timestamp 1669390400
transform 1 0 23072 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _733_
timestamp 1669390400
transform -1 0 3024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _734_
timestamp 1669390400
transform -1 0 117600 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _735_
timestamp 1669390400
transform -1 0 117600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _736_
timestamp 1669390400
transform 1 0 2352 0 1 98784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _737_
timestamp 1669390400
transform 1 0 2352 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _738_
timestamp 1669390400
transform 1 0 66752 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _739_
timestamp 1669390400
transform 1 0 111776 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _740_
timestamp 1669390400
transform 1 0 33488 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _741_
timestamp 1669390400
transform -1 0 54992 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _742_
timestamp 1669390400
transform -1 0 117600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _743_
timestamp 1669390400
transform -1 0 46480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _744_
timestamp 1669390400
transform 1 0 5488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _745_
timestamp 1669390400
transform 1 0 64288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _746_
timestamp 1669390400
transform -1 0 117600 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _747_
timestamp 1669390400
transform 1 0 76048 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _748_
timestamp 1669390400
transform 1 0 81872 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _749_
timestamp 1669390400
transform 1 0 45920 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _750_
timestamp 1669390400
transform -1 0 117600 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _751_
timestamp 1669390400
transform -1 0 45360 0 -1 103488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _752_
timestamp 1669390400
transform -1 0 117600 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _753_
timestamp 1669390400
transform 1 0 58688 0 1 89376
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _754_
timestamp 1669390400
transform 1 0 52192 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _755_
timestamp 1669390400
transform 1 0 62608 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _756_
timestamp 1669390400
transform 1 0 79856 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _757_
timestamp 1669390400
transform -1 0 117600 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _758_
timestamp 1669390400
transform -1 0 50064 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _759_
timestamp 1669390400
transform 1 0 53312 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _760_
timestamp 1669390400
transform 1 0 58128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _761_
timestamp 1669390400
transform -1 0 39984 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _762_
timestamp 1669390400
transform 1 0 53984 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _763_
timestamp 1669390400
transform 1 0 72128 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _764_
timestamp 1669390400
transform 1 0 71680 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _765_
timestamp 1669390400
transform 1 0 50512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _766_
timestamp 1669390400
transform -1 0 48832 0 -1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _767_
timestamp 1669390400
transform 1 0 89488 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _768_
timestamp 1669390400
transform -1 0 42672 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _769_
timestamp 1669390400
transform 1 0 70224 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _770_
timestamp 1669390400
transform -1 0 68320 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _771_
timestamp 1669390400
transform -1 0 69216 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 87472 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1669390400
transform -1 0 62944 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1669390400
transform 1 0 69216 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1669390400
transform -1 0 54992 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1669390400
transform 1 0 61264 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1669390400
transform -1 0 58912 0 1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1669390400
transform 1 0 57344 0 -1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1669390400
transform -1 0 66864 0 1 61152
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1669390400
transform -1 0 82768 0 1 61152
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout239
timestamp 1669390400
transform -1 0 12096 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout240
timestamp 1669390400
transform 1 0 23968 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout241
timestamp 1669390400
transform -1 0 115696 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout242
timestamp 1669390400
transform -1 0 65968 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout243
timestamp 1669390400
transform 1 0 64288 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 62384 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform -1 0 116480 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 37072 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform 1 0 49840 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform -1 0 116480 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform 1 0 41776 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform 1 0 57904 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform 1 0 1680 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform -1 0 114464 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 1680 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 116592 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform -1 0 75712 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform 1 0 56560 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform 1 0 15120 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform 1 0 10192 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform 1 0 46480 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform -1 0 56112 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input18
timestamp 1669390400
transform 1 0 1680 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input19
timestamp 1669390400
transform 1 0 1680 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input20
timestamp 1669390400
transform 1 0 1680 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input21
timestamp 1669390400
transform 1 0 1680 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input22
timestamp 1669390400
transform -1 0 116592 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input23
timestamp 1669390400
transform 1 0 43792 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input24
timestamp 1669390400
transform -1 0 116592 0 -1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input25
timestamp 1669390400
transform 1 0 21280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input26
timestamp 1669390400
transform 1 0 30800 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input27
timestamp 1669390400
transform 1 0 45136 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input28
timestamp 1669390400
transform -1 0 72464 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input29
timestamp 1669390400
transform 1 0 25200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input30
timestamp 1669390400
transform -1 0 116592 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input31
timestamp 1669390400
transform 1 0 34720 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input32
timestamp 1669390400
transform -1 0 110768 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input33
timestamp 1669390400
transform 1 0 1680 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input34
timestamp 1669390400
transform 1 0 1680 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input35
timestamp 1669390400
transform 1 0 62160 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input36
timestamp 1669390400
transform 1 0 1680 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input37
timestamp 1669390400
transform 1 0 1680 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input38
timestamp 1669390400
transform 1 0 1680 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input39
timestamp 1669390400
transform 1 0 43120 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input40 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input41
timestamp 1669390400
transform 1 0 53200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input42
timestamp 1669390400
transform 1 0 1680 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input43
timestamp 1669390400
transform -1 0 98000 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input44
timestamp 1669390400
transform 1 0 45136 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input45
timestamp 1669390400
transform 1 0 1680 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input46
timestamp 1669390400
transform -1 0 116480 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input47
timestamp 1669390400
transform -1 0 117600 0 -1 79968
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input48
timestamp 1669390400
transform -1 0 94640 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input49
timestamp 1669390400
transform 1 0 40880 0 1 116032
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input50
timestamp 1669390400
transform -1 0 116592 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input51
timestamp 1669390400
transform -1 0 83216 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input52
timestamp 1669390400
transform -1 0 116480 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input53
timestamp 1669390400
transform -1 0 93632 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input54
timestamp 1669390400
transform -1 0 109312 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input55
timestamp 1669390400
transform -1 0 116592 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input56
timestamp 1669390400
transform -1 0 75040 0 1 116032
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input57
timestamp 1669390400
transform -1 0 113232 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input58
timestamp 1669390400
transform 1 0 1680 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input59
timestamp 1669390400
transform 1 0 14896 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input60
timestamp 1669390400
transform -1 0 116592 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input61
timestamp 1669390400
transform -1 0 117600 0 -1 78400
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input62
timestamp 1669390400
transform 1 0 29680 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input63
timestamp 1669390400
transform -1 0 117152 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input64
timestamp 1669390400
transform 1 0 1680 0 1 21952
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input65
timestamp 1669390400
transform 1 0 22288 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input66
timestamp 1669390400
transform 1 0 38416 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input67
timestamp 1669390400
transform -1 0 116592 0 -1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input68
timestamp 1669390400
transform 1 0 1680 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input69
timestamp 1669390400
transform 1 0 1680 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input70
timestamp 1669390400
transform 1 0 1680 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input71
timestamp 1669390400
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input72
timestamp 1669390400
transform 1 0 1680 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input73
timestamp 1669390400
transform -1 0 116480 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input74
timestamp 1669390400
transform -1 0 71120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input75
timestamp 1669390400
transform -1 0 83888 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input76
timestamp 1669390400
transform -1 0 113456 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input77
timestamp 1669390400
transform 1 0 6160 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input78
timestamp 1669390400
transform 1 0 18256 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input79
timestamp 1669390400
transform 1 0 1680 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input80
timestamp 1669390400
transform -1 0 117152 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input81
timestamp 1669390400
transform 1 0 1680 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input82
timestamp 1669390400
transform -1 0 116480 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input83
timestamp 1669390400
transform -1 0 116592 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input84
timestamp 1669390400
transform -1 0 85792 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input85
timestamp 1669390400
transform -1 0 101472 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input86
timestamp 1669390400
transform 1 0 29008 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input87
timestamp 1669390400
transform 1 0 37744 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input88
timestamp 1669390400
transform -1 0 116480 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input89
timestamp 1669390400
transform -1 0 100016 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input90
timestamp 1669390400
transform -1 0 116480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input91
timestamp 1669390400
transform 1 0 1680 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input92
timestamp 1669390400
transform -1 0 116480 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input93
timestamp 1669390400
transform 1 0 19040 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input94
timestamp 1669390400
transform -1 0 61712 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input95
timestamp 1669390400
transform -1 0 116592 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input96
timestamp 1669390400
transform -1 0 97552 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input97
timestamp 1669390400
transform -1 0 116592 0 -1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input98
timestamp 1669390400
transform -1 0 116480 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input99
timestamp 1669390400
transform 1 0 1680 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input100
timestamp 1669390400
transform 1 0 12880 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input101
timestamp 1669390400
transform -1 0 88592 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input102
timestamp 1669390400
transform 1 0 1680 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input103
timestamp 1669390400
transform 1 0 1680 0 -1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input104
timestamp 1669390400
transform -1 0 115472 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output105 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5040 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output106
timestamp 1669390400
transform -1 0 3248 0 -1 83104
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output107
timestamp 1669390400
transform -1 0 3248 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output108
timestamp 1669390400
transform -1 0 3248 0 -1 90944
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output109
timestamp 1669390400
transform 1 0 103600 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output110
timestamp 1669390400
transform -1 0 112560 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output111
timestamp 1669390400
transform 1 0 64400 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output112
timestamp 1669390400
transform -1 0 3248 0 1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output113
timestamp 1669390400
transform 1 0 11088 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output114
timestamp 1669390400
transform -1 0 3248 0 -1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output115
timestamp 1669390400
transform 1 0 48720 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output116
timestamp 1669390400
transform -1 0 116368 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output117
timestamp 1669390400
transform 1 0 101584 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output118
timestamp 1669390400
transform 1 0 11424 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output119
timestamp 1669390400
transform -1 0 116368 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output120
timestamp 1669390400
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output121
timestamp 1669390400
transform -1 0 116368 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output122
timestamp 1669390400
transform -1 0 43568 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output123
timestamp 1669390400
transform 1 0 99680 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output124
timestamp 1669390400
transform -1 0 3248 0 1 79968
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output125
timestamp 1669390400
transform -1 0 3248 0 -1 112896
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output126
timestamp 1669390400
transform 1 0 25200 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output127
timestamp 1669390400
transform 1 0 77392 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output128
timestamp 1669390400
transform -1 0 3248 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output129
timestamp 1669390400
transform -1 0 116368 0 1 83104
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output130
timestamp 1669390400
transform -1 0 116368 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output131
timestamp 1669390400
transform -1 0 3248 0 -1 98784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output132
timestamp 1669390400
transform -1 0 3248 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output133
timestamp 1669390400
transform 1 0 68320 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output134
timestamp 1669390400
transform 1 0 113008 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output135
timestamp 1669390400
transform -1 0 116368 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output136
timestamp 1669390400
transform -1 0 3248 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output137
timestamp 1669390400
transform -1 0 116368 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output138
timestamp 1669390400
transform 1 0 57456 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output139
timestamp 1669390400
transform -1 0 116368 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output140
timestamp 1669390400
transform -1 0 116368 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output141
timestamp 1669390400
transform -1 0 116368 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output142
timestamp 1669390400
transform -1 0 3248 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output143
timestamp 1669390400
transform 1 0 114800 0 1 114464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output144
timestamp 1669390400
transform 1 0 114800 0 -1 106624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output145
timestamp 1669390400
transform 1 0 116592 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output146
timestamp 1669390400
transform -1 0 3248 0 -1 89376
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output147
timestamp 1669390400
transform -1 0 48720 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output148
timestamp 1669390400
transform 1 0 114800 0 -1 100352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output149
timestamp 1669390400
transform -1 0 15120 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output150
timestamp 1669390400
transform -1 0 103040 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output151
timestamp 1669390400
transform 1 0 78736 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output152
timestamp 1669390400
transform -1 0 9072 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output153
timestamp 1669390400
transform -1 0 83664 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output154
timestamp 1669390400
transform -1 0 56784 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output155
timestamp 1669390400
transform -1 0 42000 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output156
timestamp 1669390400
transform -1 0 3248 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output157
timestamp 1669390400
transform 1 0 88144 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output158
timestamp 1669390400
transform -1 0 56896 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output159
timestamp 1669390400
transform -1 0 52080 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output160
timestamp 1669390400
transform 1 0 85792 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output161
timestamp 1669390400
transform -1 0 90384 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output162
timestamp 1669390400
transform 1 0 76720 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output163
timestamp 1669390400
transform 1 0 113008 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output164
timestamp 1669390400
transform -1 0 112560 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output165
timestamp 1669390400
transform 1 0 114800 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output166
timestamp 1669390400
transform 1 0 100912 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output167
timestamp 1669390400
transform 1 0 114800 0 1 86240
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output168
timestamp 1669390400
transform -1 0 5040 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output169
timestamp 1669390400
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output170
timestamp 1669390400
transform -1 0 3248 0 -1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output171
timestamp 1669390400
transform 1 0 76160 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output172
timestamp 1669390400
transform -1 0 32592 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output173
timestamp 1669390400
transform -1 0 3248 0 1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output174
timestamp 1669390400
transform -1 0 35280 0 1 114464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output175
timestamp 1669390400
transform -1 0 116368 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output176
timestamp 1669390400
transform -1 0 3248 0 -1 103488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output177
timestamp 1669390400
transform -1 0 116368 0 1 67424
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output178
timestamp 1669390400
transform 1 0 59248 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output179
timestamp 1669390400
transform 1 0 53200 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output180
timestamp 1669390400
transform 1 0 63280 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output181
timestamp 1669390400
transform 1 0 114800 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output182
timestamp 1669390400
transform -1 0 116368 0 -1 114464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output183
timestamp 1669390400
transform -1 0 3248 0 1 114464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output184
timestamp 1669390400
transform 1 0 114800 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output185
timestamp 1669390400
transform -1 0 36512 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output186
timestamp 1669390400
transform 1 0 114800 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output187
timestamp 1669390400
transform -1 0 3248 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output188
timestamp 1669390400
transform 1 0 114800 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output189
timestamp 1669390400
transform 1 0 73360 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output190
timestamp 1669390400
transform 1 0 114800 0 -1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output191
timestamp 1669390400
transform 1 0 51408 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output192
timestamp 1669390400
transform -1 0 3248 0 -1 94080
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output193
timestamp 1669390400
transform 1 0 114800 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output194
timestamp 1669390400
transform -1 0 3248 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output195
timestamp 1669390400
transform -1 0 71792 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output196
timestamp 1669390400
transform -1 0 116368 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output197
timestamp 1669390400
transform -1 0 59696 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output198
timestamp 1669390400
transform -1 0 67760 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output199
timestamp 1669390400
transform -1 0 8400 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output200
timestamp 1669390400
transform 1 0 5600 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output201
timestamp 1669390400
transform 1 0 114800 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output202
timestamp 1669390400
transform -1 0 116368 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output203
timestamp 1669390400
transform 1 0 114800 0 1 84672
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output204
timestamp 1669390400
transform 1 0 114352 0 -1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output205
timestamp 1669390400
transform 1 0 47152 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output206
timestamp 1669390400
transform 1 0 114800 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output207
timestamp 1669390400
transform -1 0 3248 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output208
timestamp 1669390400
transform 1 0 114800 0 1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output209
timestamp 1669390400
transform -1 0 5264 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output210
timestamp 1669390400
transform 1 0 114800 0 -1 111328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output211
timestamp 1669390400
transform 1 0 91840 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output212
timestamp 1669390400
transform 1 0 114800 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output213
timestamp 1669390400
transform 1 0 86128 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output214
timestamp 1669390400
transform -1 0 3248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output215
timestamp 1669390400
transform -1 0 3248 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output216
timestamp 1669390400
transform 1 0 80752 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output217
timestamp 1669390400
transform -1 0 3248 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output218
timestamp 1669390400
transform 1 0 94864 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output219
timestamp 1669390400
transform -1 0 3248 0 1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output220
timestamp 1669390400
transform -1 0 3248 0 -1 105056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output221
timestamp 1669390400
transform -1 0 33040 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output222
timestamp 1669390400
transform -1 0 3248 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output223
timestamp 1669390400
transform -1 0 26544 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output224
timestamp 1669390400
transform -1 0 11088 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output225
timestamp 1669390400
transform -1 0 64176 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output226
timestamp 1669390400
transform -1 0 36624 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output227
timestamp 1669390400
transform 1 0 64624 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output228
timestamp 1669390400
transform 1 0 84000 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output229
timestamp 1669390400
transform -1 0 116368 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output230
timestamp 1669390400
transform -1 0 3248 0 1 78400
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output231
timestamp 1669390400
transform 1 0 114800 0 1 92512
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output232
timestamp 1669390400
transform -1 0 27888 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output233
timestamp 1669390400
transform 1 0 46480 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output234
timestamp 1669390400
transform -1 0 3248 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output235
timestamp 1669390400
transform -1 0 116368 0 1 89376
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output236
timestamp 1669390400
transform 1 0 73248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output237
timestamp 1669390400
transform -1 0 80304 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output238
timestamp 1669390400
transform 1 0 78064 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_244 gf180mcu-pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2128 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_245
timestamp 1669390400
transform 1 0 117824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_246
timestamp 1669390400
transform -1 0 80528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_247
timestamp 1669390400
transform 1 0 117824 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_248
timestamp 1669390400
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_249
timestamp 1669390400
transform 1 0 117824 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_250
timestamp 1669390400
transform 1 0 117824 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_251
timestamp 1669390400
transform -1 0 2128 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_252
timestamp 1669390400
transform -1 0 2128 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_253
timestamp 1669390400
transform -1 0 37520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_254
timestamp 1669390400
transform 1 0 117824 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_255
timestamp 1669390400
transform 1 0 117824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_256
timestamp 1669390400
transform 1 0 117824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_257
timestamp 1669390400
transform 1 0 117824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_258
timestamp 1669390400
transform -1 0 2128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_259
timestamp 1669390400
transform -1 0 2128 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_260
timestamp 1669390400
transform -1 0 2128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_261
timestamp 1669390400
transform 1 0 117824 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_262
timestamp 1669390400
transform -1 0 50288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_263
timestamp 1669390400
transform -1 0 19376 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_264
timestamp 1669390400
transform -1 0 110096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_265
timestamp 1669390400
transform -1 0 2128 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_266
timestamp 1669390400
transform -1 0 28000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_267
timestamp 1669390400
transform -1 0 109424 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_268
timestamp 1669390400
transform -1 0 69888 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_269
timestamp 1669390400
transform -1 0 42224 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_270
timestamp 1669390400
transform -1 0 5040 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_271
timestamp 1669390400
transform -1 0 87248 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_272
timestamp 1669390400
transform -1 0 94640 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_273
timestamp 1669390400
transform -1 0 51632 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_274
timestamp 1669390400
transform -1 0 2128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_275
timestamp 1669390400
transform 1 0 117824 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_276
timestamp 1669390400
transform 1 0 117824 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_277
timestamp 1669390400
transform 1 0 117824 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_278
timestamp 1669390400
transform -1 0 2128 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_279
timestamp 1669390400
transform -1 0 98224 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_280
timestamp 1669390400
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_281
timestamp 1669390400
transform -1 0 105840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_282
timestamp 1669390400
transform -1 0 2128 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_283
timestamp 1669390400
transform -1 0 44352 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_284
timestamp 1669390400
transform -1 0 76608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_285
timestamp 1669390400
transform 1 0 117824 0 1 56448
box -86 -86 534 870
<< labels >>
flabel metal3 s 200 41608 800 41832 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 200 55048 800 55272 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 200 49672 800 49896 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 115528 119200 115752 119800 0 FreeSans 896 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 200 42280 800 42504 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 65800 119200 66024 119800 0 FreeSans 896 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal3 s 119200 22792 119800 23016 0 FreeSans 896 0 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 34216 200 34440 800 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 26824 119200 27048 119800 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal3 s 200 53032 800 53256 0 FreeSans 896 0 0 0 io_in[18]
port 9 nsew signal input
flabel metal3 s 119200 119560 119800 119784 0 FreeSans 896 0 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 96040 119200 96264 119800 0 FreeSans 896 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 69160 119200 69384 119800 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 113512 119200 113736 119800 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 1960 119200 2184 119800 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 16072 200 16296 800 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 14728 119200 14952 119800 0 FreeSans 896 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 19432 119200 19656 119800 0 FreeSans 896 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 119200 12712 119800 12936 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 200 28840 800 29064 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 4648 119200 4872 119800 0 FreeSans 896 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 119200 116872 119800 117096 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 200 12040 800 12264 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 83944 200 84168 800 0 FreeSans 896 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 17416 119200 17640 119800 0 FreeSans 896 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 71176 200 71400 800 0 FreeSans 896 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 200 117544 800 117768 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 107464 119200 107688 119800 0 FreeSans 896 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 25480 119200 25704 119800 0 FreeSans 896 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 200 30856 800 31080 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 119200 19432 119800 19656 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 200 50344 800 50568 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 107464 200 107688 800 0 FreeSans 896 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 200 116872 800 117096 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 200 27496 800 27720 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 119200 31528 119800 31752 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 116872 200 117096 800 0 FreeSans 896 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 102088 119200 102312 119800 0 FreeSans 896 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 3304 119200 3528 119800 0 FreeSans 896 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 200 81928 800 82152 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 200 75208 800 75432 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 200 89992 800 90216 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 102760 200 102984 800 0 FreeSans 896 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 117544 200 117768 800 0 FreeSans 896 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 63784 119200 64008 119800 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal3 s 200 69160 800 69384 0 FreeSans 896 0 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 11368 119200 11592 119800 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal3 s 200 94696 800 94920 0 FreeSans 896 0 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 48328 200 48552 800 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 119200 9352 119800 9576 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 101416 200 101640 800 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 11368 200 11592 800 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal3 s 119200 30184 119800 30408 0 FreeSans 896 0 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal3 s 200 11368 800 11592 0 FreeSans 896 0 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 119200 26824 119800 27048 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 42280 200 42504 800 0 FreeSans 896 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 99400 200 99624 800 0 FreeSans 896 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 200 79912 800 80136 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 200 112168 800 112392 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 24136 119200 24360 119800 0 FreeSans 896 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 77224 200 77448 800 0 FreeSans 896 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 200 3976 800 4200 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 119200 83272 119800 83496 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 119200 18760 119800 18984 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 200 98056 800 98280 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 200 46312 800 46536 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 67144 119200 67368 119800 0 FreeSans 896 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 112168 200 112392 800 0 FreeSans 896 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 200 100744 800 100968 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 119200 40264 119800 40488 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s -56 119200 168 119800 0 FreeSans 896 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 119200 115528 119800 115752 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 57736 119200 57960 119800 0 FreeSans 896 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 119200 6664 119800 6888 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 119200 48328 119800 48552 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 119200 47656 119800 47880 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 200 22792 800 23016 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 116872 119200 117096 119800 0 FreeSans 896 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 119200 105448 119800 105672 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 119200 118216 119800 118440 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 200 88648 800 88872 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 46984 200 47208 800 0 FreeSans 896 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal3 s 119200 99400 119800 99624 0 FreeSans 896 0 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 13384 200 13608 800 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 100744 200 100968 800 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 78568 200 78792 800 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 8008 200 8232 800 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 81928 200 82152 800 0 FreeSans 896 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 54376 200 54600 800 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 40264 200 40488 800 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal3 s 200 16072 800 16296 0 FreeSans 896 0 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 87976 119200 88200 119800 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 55720 119200 55944 119800 0 FreeSans 896 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 50344 200 50568 800 0 FreeSans 896 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 84616 119200 84840 119800 0 FreeSans 896 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 88648 200 88872 800 0 FreeSans 896 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 76552 119200 76776 119800 0 FreeSans 896 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 113512 200 113736 800 0 FreeSans 896 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 110152 119200 110376 119800 0 FreeSans 896 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 119200 25480 119800 25704 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 100744 119200 100968 119800 0 FreeSans 896 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 119200 38248 119800 38472 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 79912 200 80136 800 0 FreeSans 896 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 119200 77896 119800 78120 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 28840 200 29064 800 0 FreeSans 896 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 119200 112168 119800 112392 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 119200 111496 119800 111720 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 119200 85960 119800 86184 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 200 3304 800 3528 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 200 5320 800 5544 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 200 67816 800 68040 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 75208 119200 75432 119800 0 FreeSans 896 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 30856 200 31080 800 0 FreeSans 896 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 200 61096 800 61320 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal3 s 200 83944 800 84168 0 FreeSans 896 0 0 0 irq[0]
port 114 nsew signal tristate
flabel metal3 s 200 48328 800 48552 0 FreeSans 896 0 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 36904 200 37128 800 0 FreeSans 896 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 48328 119200 48552 119800 0 FreeSans 896 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 112168 119200 112392 119800 0 FreeSans 896 90 0 0 la_data_in[10]
port 118 nsew signal input
flabel metal2 s 56392 200 56616 800 0 FreeSans 896 90 0 0 la_data_in[11]
port 119 nsew signal input
flabel metal3 s 200 72520 800 72744 0 FreeSans 896 0 0 0 la_data_in[12]
port 120 nsew signal input
flabel metal3 s 119200 17416 119800 17640 0 FreeSans 896 0 0 0 la_data_in[13]
port 121 nsew signal input
flabel metal3 s 119200 43624 119800 43848 0 FreeSans 896 0 0 0 la_data_in[14]
port 122 nsew signal input
flabel metal3 s 200 83272 800 83496 0 FreeSans 896 0 0 0 la_data_in[15]
port 123 nsew signal input
flabel metal2 s 27496 119200 27720 119800 0 FreeSans 896 90 0 0 la_data_in[16]
port 124 nsew signal input
flabel metal3 s 119200 24136 119800 24360 0 FreeSans 896 0 0 0 la_data_in[17]
port 125 nsew signal input
flabel metal3 s 119200 90664 119800 90888 0 FreeSans 896 0 0 0 la_data_in[18]
port 126 nsew signal input
flabel metal3 s 119200 53032 119800 53256 0 FreeSans 896 0 0 0 la_data_in[19]
port 127 nsew signal input
flabel metal2 s 91336 119200 91560 119800 0 FreeSans 896 90 0 0 la_data_in[1]
port 128 nsew signal input
flabel metal2 s 61096 119200 61320 119800 0 FreeSans 896 90 0 0 la_data_in[20]
port 129 nsew signal input
flabel metal3 s 200 19432 800 19656 0 FreeSans 896 0 0 0 la_data_in[21]
port 130 nsew signal input
flabel metal2 s 73864 119200 74088 119800 0 FreeSans 896 90 0 0 la_data_in[22]
port 131 nsew signal input
flabel metal3 s 200 108808 800 109032 0 FreeSans 896 0 0 0 la_data_in[23]
port 132 nsew signal input
flabel metal2 s 52360 119200 52584 119800 0 FreeSans 896 90 0 0 la_data_in[24]
port 133 nsew signal input
flabel metal3 s 119200 28840 119800 29064 0 FreeSans 896 0 0 0 la_data_in[25]
port 134 nsew signal input
flabel metal2 s 38920 200 39144 800 0 FreeSans 896 90 0 0 la_data_in[26]
port 135 nsew signal input
flabel metal3 s 200 8680 800 8904 0 FreeSans 896 0 0 0 la_data_in[27]
port 136 nsew signal input
flabel metal3 s 200 43624 800 43848 0 FreeSans 896 0 0 0 la_data_in[28]
port 137 nsew signal input
flabel metal3 s 200 91336 800 91560 0 FreeSans 896 0 0 0 la_data_in[29]
port 138 nsew signal input
flabel metal3 s 200 80584 800 80808 0 FreeSans 896 0 0 0 la_data_in[2]
port 139 nsew signal input
flabel metal2 s 9352 119200 9576 119800 0 FreeSans 896 90 0 0 la_data_in[30]
port 140 nsew signal input
flabel metal3 s 200 106120 800 106344 0 FreeSans 896 0 0 0 la_data_in[31]
port 141 nsew signal input
flabel metal2 s 60424 119200 60648 119800 0 FreeSans 896 90 0 0 la_data_in[32]
port 142 nsew signal input
flabel metal3 s 119200 102088 119800 102312 0 FreeSans 896 0 0 0 la_data_in[33]
port 143 nsew signal input
flabel metal2 s 36904 119200 37128 119800 0 FreeSans 896 90 0 0 la_data_in[34]
port 144 nsew signal input
flabel metal2 s 49672 119200 49896 119800 0 FreeSans 896 90 0 0 la_data_in[35]
port 145 nsew signal input
flabel metal3 s 119200 65128 119800 65352 0 FreeSans 896 0 0 0 la_data_in[36]
port 146 nsew signal input
flabel metal2 s 41608 200 41832 800 0 FreeSans 896 90 0 0 la_data_in[37]
port 147 nsew signal input
flabel metal2 s 57736 200 57960 800 0 FreeSans 896 90 0 0 la_data_in[38]
port 148 nsew signal input
flabel metal3 s 200 40264 800 40488 0 FreeSans 896 0 0 0 la_data_in[39]
port 149 nsew signal input
flabel metal3 s 119200 73864 119800 74088 0 FreeSans 896 0 0 0 la_data_in[3]
port 150 nsew signal input
flabel metal3 s 119200 1288 119800 1512 0 FreeSans 896 0 0 0 la_data_in[40]
port 151 nsew signal input
flabel metal3 s 200 113512 800 113736 0 FreeSans 896 0 0 0 la_data_in[41]
port 152 nsew signal input
flabel metal3 s 119200 86632 119800 86856 0 FreeSans 896 0 0 0 la_data_in[42]
port 153 nsew signal input
flabel metal2 s 73864 200 74088 800 0 FreeSans 896 90 0 0 la_data_in[43]
port 154 nsew signal input
flabel metal2 s 56392 119200 56616 119800 0 FreeSans 896 90 0 0 la_data_in[44]
port 155 nsew signal input
flabel metal2 s 16072 119200 16296 119800 0 FreeSans 896 90 0 0 la_data_in[45]
port 156 nsew signal input
flabel metal2 s 10024 119200 10248 119800 0 FreeSans 896 90 0 0 la_data_in[46]
port 157 nsew signal input
flabel metal2 s 47656 119200 47880 119800 0 FreeSans 896 90 0 0 la_data_in[47]
port 158 nsew signal input
flabel metal2 s 55048 200 55272 800 0 FreeSans 896 90 0 0 la_data_in[48]
port 159 nsew signal input
flabel metal3 s 200 62440 800 62664 0 FreeSans 896 0 0 0 la_data_in[49]
port 160 nsew signal input
flabel metal2 s 98728 119200 98952 119800 0 FreeSans 896 90 0 0 la_data_in[4]
port 161 nsew signal input
flabel metal3 s 200 36904 800 37128 0 FreeSans 896 0 0 0 la_data_in[50]
port 162 nsew signal input
flabel metal3 s 200 32200 800 32424 0 FreeSans 896 0 0 0 la_data_in[51]
port 163 nsew signal input
flabel metal3 s 200 35560 800 35784 0 FreeSans 896 0 0 0 la_data_in[52]
port 164 nsew signal input
flabel metal3 s 119200 3304 119800 3528 0 FreeSans 896 0 0 0 la_data_in[53]
port 165 nsew signal input
flabel metal2 s 43624 200 43848 800 0 FreeSans 896 90 0 0 la_data_in[54]
port 166 nsew signal input
flabel metal3 s 119200 108808 119800 109032 0 FreeSans 896 0 0 0 la_data_in[55]
port 167 nsew signal input
flabel metal2 s 20776 200 21000 800 0 FreeSans 896 90 0 0 la_data_in[56]
port 168 nsew signal input
flabel metal2 s 31528 119200 31752 119800 0 FreeSans 896 90 0 0 la_data_in[57]
port 169 nsew signal input
flabel metal2 s 44968 119200 45192 119800 0 FreeSans 896 90 0 0 la_data_in[58]
port 170 nsew signal input
flabel metal2 s 70504 200 70728 800 0 FreeSans 896 90 0 0 la_data_in[59]
port 171 nsew signal input
flabel metal3 s 200 616 800 840 0 FreeSans 896 0 0 0 la_data_in[5]
port 172 nsew signal input
flabel metal2 s 24136 200 24360 800 0 FreeSans 896 90 0 0 la_data_in[60]
port 173 nsew signal input
flabel metal3 s 119200 42952 119800 43176 0 FreeSans 896 0 0 0 la_data_in[61]
port 174 nsew signal input
flabel metal2 s 35560 119200 35784 119800 0 FreeSans 896 90 0 0 la_data_in[62]
port 175 nsew signal input
flabel metal2 s 108808 119200 109032 119800 0 FreeSans 896 90 0 0 la_data_in[63]
port 176 nsew signal input
flabel metal2 s 104104 119200 104328 119800 0 FreeSans 896 90 0 0 la_data_in[6]
port 177 nsew signal input
flabel metal3 s 119200 63784 119800 64008 0 FreeSans 896 0 0 0 la_data_in[7]
port 178 nsew signal input
flabel metal2 s 85288 200 85512 800 0 FreeSans 896 90 0 0 la_data_in[8]
port 179 nsew signal input
flabel metal3 s 200 86632 800 86856 0 FreeSans 896 0 0 0 la_data_in[9]
port 180 nsew signal input
flabel metal2 s 33544 119200 33768 119800 0 FreeSans 896 90 0 0 la_data_out[0]
port 181 nsew signal tristate
flabel metal3 s 119200 49672 119800 49896 0 FreeSans 896 0 0 0 la_data_out[10]
port 182 nsew signal tristate
flabel metal3 s 200 102760 800 102984 0 FreeSans 896 0 0 0 la_data_out[11]
port 183 nsew signal tristate
flabel metal3 s 119200 65800 119800 66024 0 FreeSans 896 0 0 0 la_data_out[12]
port 184 nsew signal tristate
flabel metal2 s 59080 119200 59304 119800 0 FreeSans 896 90 0 0 la_data_out[13]
port 185 nsew signal tristate
flabel metal2 s 53032 119200 53256 119800 0 FreeSans 896 90 0 0 la_data_out[14]
port 186 nsew signal tristate
flabel metal2 s 63112 200 63336 800 0 FreeSans 896 90 0 0 la_data_out[15]
port 187 nsew signal tristate
flabel metal3 s 119200 55720 119800 55944 0 FreeSans 896 0 0 0 la_data_out[16]
port 188 nsew signal tristate
flabel metal2 s 118216 119200 118440 119800 0 FreeSans 896 90 0 0 la_data_out[17]
port 189 nsew signal tristate
flabel metal3 s 200 118888 800 119112 0 FreeSans 896 0 0 0 la_data_out[18]
port 190 nsew signal tristate
flabel metal3 s 119200 75208 119800 75432 0 FreeSans 896 0 0 0 la_data_out[19]
port 191 nsew signal tristate
flabel metal2 s 35560 200 35784 800 0 FreeSans 896 90 0 0 la_data_out[1]
port 192 nsew signal tristate
flabel metal3 s 119200 34888 119800 35112 0 FreeSans 896 0 0 0 la_data_out[20]
port 193 nsew signal tristate
flabel metal3 s 200 20776 800 21000 0 FreeSans 896 0 0 0 la_data_out[21]
port 194 nsew signal tristate
flabel metal3 s 119200 14728 119800 14952 0 FreeSans 896 0 0 0 la_data_out[22]
port 195 nsew signal tristate
flabel metal2 s 73192 119200 73416 119800 0 FreeSans 896 90 0 0 la_data_out[23]
port 196 nsew signal tristate
flabel metal3 s 119200 94696 119800 94920 0 FreeSans 896 0 0 0 la_data_out[24]
port 197 nsew signal tristate
flabel metal2 s 51688 200 51912 800 0 FreeSans 896 90 0 0 la_data_out[25]
port 198 nsew signal tristate
flabel metal3 s 200 93352 800 93576 0 FreeSans 896 0 0 0 la_data_out[26]
port 199 nsew signal tristate
flabel metal3 s 119200 54376 119800 54600 0 FreeSans 896 0 0 0 la_data_out[27]
port 200 nsew signal tristate
flabel metal3 s 200 44968 800 45192 0 FreeSans 896 0 0 0 la_data_out[28]
port 201 nsew signal tristate
flabel metal2 s 70504 119200 70728 119800 0 FreeSans 896 90 0 0 la_data_out[29]
port 202 nsew signal tristate
flabel metal3 s 119200 22120 119800 22344 0 FreeSans 896 0 0 0 la_data_out[2]
port 203 nsew signal tristate
flabel metal2 s 58408 200 58632 800 0 FreeSans 896 90 0 0 la_data_out[30]
port 204 nsew signal tristate
flabel metal2 s 65128 119200 65352 119800 0 FreeSans 896 90 0 0 la_data_out[31]
port 205 nsew signal tristate
flabel metal3 s 119200 96040 119800 96264 0 FreeSans 896 0 0 0 la_data_out[32]
port 206 nsew signal tristate
flabel metal3 s 119200 46312 119800 46536 0 FreeSans 896 0 0 0 la_data_out[33]
port 207 nsew signal tristate
flabel metal3 s 119200 1960 119800 2184 0 FreeSans 896 0 0 0 la_data_out[34]
port 208 nsew signal tristate
flabel metal3 s 119200 16072 119800 16296 0 FreeSans 896 0 0 0 la_data_out[35]
port 209 nsew signal tristate
flabel metal3 s 200 6664 800 6888 0 FreeSans 896 0 0 0 la_data_out[36]
port 210 nsew signal tristate
flabel metal3 s 200 107464 800 107688 0 FreeSans 896 0 0 0 la_data_out[37]
port 211 nsew signal tristate
flabel metal3 s 200 54376 800 54600 0 FreeSans 896 0 0 0 la_data_out[38]
port 212 nsew signal tristate
flabel metal3 s 119200 100744 119800 100968 0 FreeSans 896 0 0 0 la_data_out[39]
port 213 nsew signal tristate
flabel metal2 s 6664 200 6888 800 0 FreeSans 896 90 0 0 la_data_out[3]
port 214 nsew signal tristate
flabel metal2 s 49672 200 49896 800 0 FreeSans 896 90 0 0 la_data_out[40]
port 215 nsew signal tristate
flabel metal2 s 18760 119200 18984 119800 0 FreeSans 896 90 0 0 la_data_out[41]
port 216 nsew signal tristate
flabel metal2 s 109480 200 109704 800 0 FreeSans 896 90 0 0 la_data_out[42]
port 217 nsew signal tristate
flabel metal3 s 200 85288 800 85512 0 FreeSans 896 0 0 0 la_data_out[43]
port 218 nsew signal tristate
flabel metal2 s 27496 200 27720 800 0 FreeSans 896 90 0 0 la_data_out[44]
port 219 nsew signal tristate
flabel metal2 s 108808 200 109032 800 0 FreeSans 896 90 0 0 la_data_out[45]
port 220 nsew signal tristate
flabel metal2 s 68488 119200 68712 119800 0 FreeSans 896 90 0 0 la_data_out[46]
port 221 nsew signal tristate
flabel metal2 s 41608 119200 41832 119800 0 FreeSans 896 90 0 0 la_data_out[47]
port 222 nsew signal tristate
flabel metal3 s 200 115528 800 115752 0 FreeSans 896 0 0 0 la_data_out[48]
port 223 nsew signal tristate
flabel metal2 s 86632 119200 86856 119800 0 FreeSans 896 90 0 0 la_data_out[49]
port 224 nsew signal tristate
flabel metal3 s 200 1960 800 2184 0 FreeSans 896 0 0 0 la_data_out[4]
port 225 nsew signal tristate
flabel metal2 s 94024 119200 94248 119800 0 FreeSans 896 90 0 0 la_data_out[50]
port 226 nsew signal tristate
flabel metal2 s 51016 119200 51240 119800 0 FreeSans 896 90 0 0 la_data_out[51]
port 227 nsew signal tristate
flabel metal3 s 200 16744 800 16968 0 FreeSans 896 0 0 0 la_data_out[52]
port 228 nsew signal tristate
flabel metal3 s 119200 70504 119800 70728 0 FreeSans 896 0 0 0 la_data_out[53]
port 229 nsew signal tristate
flabel metal3 s 119200 81928 119800 82152 0 FreeSans 896 0 0 0 la_data_out[54]
port 230 nsew signal tristate
flabel metal3 s 119200 106792 119800 107016 0 FreeSans 896 0 0 0 la_data_out[55]
port 231 nsew signal tristate
flabel metal3 s 200 109480 800 109704 0 FreeSans 896 0 0 0 la_data_out[56]
port 232 nsew signal tristate
flabel metal2 s 97384 119200 97608 119800 0 FreeSans 896 90 0 0 la_data_out[57]
port 233 nsew signal tristate
flabel metal2 s 32200 200 32424 800 0 FreeSans 896 90 0 0 la_data_out[58]
port 234 nsew signal tristate
flabel metal2 s 104104 200 104328 800 0 FreeSans 896 90 0 0 la_data_out[59]
port 235 nsew signal tristate
flabel metal3 s 119200 8008 119800 8232 0 FreeSans 896 0 0 0 la_data_out[5]
port 236 nsew signal tristate
flabel metal3 s 200 18088 800 18312 0 FreeSans 896 0 0 0 la_data_out[60]
port 237 nsew signal tristate
flabel metal2 s 42952 119200 43176 119800 0 FreeSans 896 90 0 0 la_data_out[61]
port 238 nsew signal tristate
flabel metal2 s 75208 200 75432 800 0 FreeSans 896 90 0 0 la_data_out[62]
port 239 nsew signal tristate
flabel metal3 s 119200 56392 119800 56616 0 FreeSans 896 0 0 0 la_data_out[63]
port 240 nsew signal tristate
flabel metal3 s 119200 44968 119800 45192 0 FreeSans 896 0 0 0 la_data_out[6]
port 241 nsew signal tristate
flabel metal3 s 119200 84616 119800 84840 0 FreeSans 896 0 0 0 la_data_out[7]
port 242 nsew signal tristate
flabel metal3 s 119200 67144 119800 67368 0 FreeSans 896 0 0 0 la_data_out[8]
port 243 nsew signal tristate
flabel metal2 s 46312 119200 46536 119800 0 FreeSans 896 90 0 0 la_data_out[9]
port 244 nsew signal tristate
flabel metal3 s 200 96040 800 96264 0 FreeSans 896 0 0 0 la_oenb[0]
port 245 nsew signal input
flabel metal2 s 87976 200 88200 800 0 FreeSans 896 90 0 0 la_oenb[10]
port 246 nsew signal input
flabel metal2 s 105448 200 105672 800 0 FreeSans 896 90 0 0 la_oenb[11]
port 247 nsew signal input
flabel metal2 s 16744 200 16968 800 0 FreeSans 896 90 0 0 la_oenb[12]
port 248 nsew signal input
flabel metal3 s 200 14728 800 14952 0 FreeSans 896 0 0 0 la_oenb[13]
port 249 nsew signal input
flabel metal2 s 8008 119200 8232 119800 0 FreeSans 896 90 0 0 la_oenb[14]
port 250 nsew signal input
flabel metal3 s 119200 10024 119800 10248 0 FreeSans 896 0 0 0 la_oenb[15]
port 251 nsew signal input
flabel metal2 s 22792 119200 23016 119800 0 FreeSans 896 90 0 0 la_oenb[16]
port 252 nsew signal input
flabel metal3 s 200 105448 800 105672 0 FreeSans 896 0 0 0 la_oenb[17]
port 253 nsew signal input
flabel metal2 s 105448 119200 105672 119800 0 FreeSans 896 90 0 0 la_oenb[18]
port 254 nsew signal input
flabel metal2 s 89320 119200 89544 119800 0 FreeSans 896 90 0 0 la_oenb[19]
port 255 nsew signal input
flabel metal2 s 33544 200 33768 800 0 FreeSans 896 90 0 0 la_oenb[1]
port 256 nsew signal input
flabel metal3 s 200 67144 800 67368 0 FreeSans 896 0 0 0 la_oenb[20]
port 257 nsew signal input
flabel metal2 s 106120 200 106344 800 0 FreeSans 896 90 0 0 la_oenb[21]
port 258 nsew signal input
flabel metal3 s 200 64456 800 64680 0 FreeSans 896 0 0 0 la_oenb[22]
port 259 nsew signal input
flabel metal2 s 21448 200 21672 800 0 FreeSans 896 90 0 0 la_oenb[23]
port 260 nsew signal input
flabel metal3 s 200 73864 800 74088 0 FreeSans 896 0 0 0 la_oenb[24]
port 261 nsew signal input
flabel metal3 s 119200 113512 119800 113736 0 FreeSans 896 0 0 0 la_oenb[25]
port 262 nsew signal input
flabel metal2 s 119560 119200 119784 119800 0 FreeSans 896 90 0 0 la_oenb[26]
port 263 nsew signal input
flabel metal3 s 119200 102760 119800 102984 0 FreeSans 896 0 0 0 la_oenb[27]
port 264 nsew signal input
flabel metal3 s 119200 98728 119800 98952 0 FreeSans 896 0 0 0 la_oenb[28]
port 265 nsew signal input
flabel metal3 s 119200 97384 119800 97608 0 FreeSans 896 0 0 0 la_oenb[29]
port 266 nsew signal input
flabel metal2 s 61096 200 61320 800 0 FreeSans 896 90 0 0 la_oenb[2]
port 267 nsew signal input
flabel metal2 s 20776 119200 21000 119800 0 FreeSans 896 90 0 0 la_oenb[30]
port 268 nsew signal input
flabel metal2 s 3304 200 3528 800 0 FreeSans 896 90 0 0 la_oenb[31]
port 269 nsew signal input
flabel metal2 s 616 200 840 800 0 FreeSans 896 90 0 0 la_oenb[32]
port 270 nsew signal input
flabel metal2 s 1288 119200 1512 119800 0 FreeSans 896 90 0 0 la_oenb[33]
port 271 nsew signal input
flabel metal2 s 62440 200 62664 800 0 FreeSans 896 90 0 0 la_oenb[34]
port 272 nsew signal input
flabel metal3 s 200 51688 800 51912 0 FreeSans 896 0 0 0 la_oenb[35]
port 273 nsew signal input
flabel metal3 s 200 65800 800 66024 0 FreeSans 896 0 0 0 la_oenb[36]
port 274 nsew signal input
flabel metal3 s 200 34216 800 34440 0 FreeSans 896 0 0 0 la_oenb[37]
port 275 nsew signal input
flabel metal2 s 43624 119200 43848 119800 0 FreeSans 896 90 0 0 la_oenb[38]
port 276 nsew signal input
flabel metal3 s 200 75880 800 76104 0 FreeSans 896 0 0 0 la_oenb[39]
port 277 nsew signal input
flabel metal2 s 22792 200 23016 800 0 FreeSans 896 90 0 0 la_oenb[3]
port 278 nsew signal input
flabel metal2 s 53032 200 53256 800 0 FreeSans 896 90 0 0 la_oenb[40]
port 279 nsew signal input
flabel metal3 s 200 59752 800 59976 0 FreeSans 896 0 0 0 la_oenb[41]
port 280 nsew signal input
flabel metal2 s 96040 200 96264 800 0 FreeSans 896 90 0 0 la_oenb[42]
port 281 nsew signal input
flabel metal2 s 44968 200 45192 800 0 FreeSans 896 90 0 0 la_oenb[43]
port 282 nsew signal input
flabel metal3 s 200 87976 800 88200 0 FreeSans 896 0 0 0 la_oenb[44]
port 283 nsew signal input
flabel metal3 s 119200 57736 119800 57960 0 FreeSans 896 0 0 0 la_oenb[45]
port 284 nsew signal input
flabel metal3 s 119200 79912 119800 80136 0 FreeSans 896 0 0 0 la_oenb[46]
port 285 nsew signal input
flabel metal2 s 92680 200 92904 800 0 FreeSans 896 90 0 0 la_oenb[47]
port 286 nsew signal input
flabel metal2 s 39592 119200 39816 119800 0 FreeSans 896 90 0 0 la_oenb[48]
port 287 nsew signal input
flabel metal2 s 118888 200 119112 800 0 FreeSans 896 90 0 0 la_oenb[49]
port 288 nsew signal input
flabel metal3 s 119200 76552 119800 76776 0 FreeSans 896 0 0 0 la_oenb[4]
port 289 nsew signal input
flabel metal2 s 81256 119200 81480 119800 0 FreeSans 896 90 0 0 la_oenb[50]
port 290 nsew signal input
flabel metal3 s 119200 61096 119800 61320 0 FreeSans 896 0 0 0 la_oenb[51]
port 291 nsew signal input
flabel metal2 s 91336 200 91560 800 0 FreeSans 896 90 0 0 la_oenb[52]
port 292 nsew signal input
flabel metal2 s 106792 119200 107016 119800 0 FreeSans 896 90 0 0 la_oenb[53]
port 293 nsew signal input
flabel metal3 s 119200 11368 119800 11592 0 FreeSans 896 0 0 0 la_oenb[54]
port 294 nsew signal input
flabel metal2 s 71848 119200 72072 119800 0 FreeSans 896 90 0 0 la_oenb[55]
port 295 nsew signal input
flabel metal2 s 110824 200 111048 800 0 FreeSans 896 90 0 0 la_oenb[56]
port 296 nsew signal input
flabel metal3 s 200 58408 800 58632 0 FreeSans 896 0 0 0 la_oenb[57]
port 297 nsew signal input
flabel metal2 s 14728 200 14952 800 0 FreeSans 896 90 0 0 la_oenb[58]
port 298 nsew signal input
flabel metal3 s 119200 60424 119800 60648 0 FreeSans 896 0 0 0 la_oenb[59]
port 299 nsew signal input
flabel metal3 s 200 114184 800 114408 0 FreeSans 896 0 0 0 la_oenb[5]
port 300 nsew signal input
flabel metal3 s 119200 78568 119800 78792 0 FreeSans 896 0 0 0 la_oenb[60]
port 301 nsew signal input
flabel metal2 s 29512 200 29736 800 0 FreeSans 896 90 0 0 la_oenb[61]
port 302 nsew signal input
flabel metal2 s 114184 200 114408 800 0 FreeSans 896 90 0 0 la_oenb[62]
port 303 nsew signal input
flabel metal3 s 200 21448 800 21672 0 FreeSans 896 0 0 0 la_oenb[63]
port 304 nsew signal input
flabel metal2 s 102760 119200 102984 119800 0 FreeSans 896 90 0 0 la_oenb[6]
port 305 nsew signal input
flabel metal3 s 119200 91336 119800 91560 0 FreeSans 896 0 0 0 la_oenb[7]
port 306 nsew signal input
flabel metal2 s 30184 119200 30408 119800 0 FreeSans 896 90 0 0 la_oenb[8]
port 307 nsew signal input
flabel metal3 s 200 77224 800 77448 0 FreeSans 896 0 0 0 la_oenb[9]
port 308 nsew signal input
flabel metal4 s 4448 3076 4768 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 35168 3076 35488 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 65888 3076 66208 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 96608 3076 96928 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 19808 3076 20128 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal3 s 119200 20776 119800 21000 0 FreeSans 896 0 0 0 wb_clk_i
port 311 nsew signal input
flabel metal2 s 22120 119200 22344 119800 0 FreeSans 896 90 0 0 wb_rst_i
port 312 nsew signal input
flabel metal3 s 119200 41608 119800 41832 0 FreeSans 896 0 0 0 wbs_ack_o
port 313 nsew signal tristate
flabel metal2 s 79912 119200 80136 119800 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 314 nsew signal input
flabel metal2 s 54376 119200 54600 119800 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 315 nsew signal input
flabel metal2 s 6664 119200 6888 119800 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 316 nsew signal input
flabel metal2 s 10024 200 10248 800 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 317 nsew signal input
flabel metal2 s 67144 200 67368 800 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 318 nsew signal input
flabel metal3 s 119200 87976 119800 88200 0 FreeSans 896 0 0 0 wbs_adr_i[14]
port 319 nsew signal input
flabel metal3 s 119200 81256 119800 81480 0 FreeSans 896 0 0 0 wbs_adr_i[15]
port 320 nsew signal input
flabel metal2 s 75880 200 76104 800 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 321 nsew signal input
flabel metal3 s 119200 71848 119800 72072 0 FreeSans 896 0 0 0 wbs_adr_i[17]
port 322 nsew signal input
flabel metal3 s 119200 36904 119800 37128 0 FreeSans 896 0 0 0 wbs_adr_i[18]
port 323 nsew signal input
flabel metal2 s 115528 200 115752 800 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 324 nsew signal input
flabel metal3 s 200 8008 800 8232 0 FreeSans 896 0 0 0 wbs_adr_i[1]
port 325 nsew signal input
flabel metal3 s 200 70504 800 70728 0 FreeSans 896 0 0 0 wbs_adr_i[20]
port 326 nsew signal input
flabel metal2 s 67816 200 68040 800 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 327 nsew signal input
flabel metal2 s 96712 200 96936 800 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 328 nsew signal input
flabel metal3 s 119200 27496 119800 27720 0 FreeSans 896 0 0 0 wbs_adr_i[23]
port 329 nsew signal input
flabel metal2 s 14056 119200 14280 119800 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 330 nsew signal input
flabel metal2 s 65800 200 66024 800 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 331 nsew signal input
flabel metal2 s 12040 200 12264 800 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 332 nsew signal input
flabel metal2 s 40264 119200 40488 119800 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 333 nsew signal input
flabel metal3 s 119200 69160 119800 69384 0 FreeSans 896 0 0 0 wbs_adr_i[28]
port 334 nsew signal input
flabel metal3 s 119200 114856 119800 115080 0 FreeSans 896 0 0 0 wbs_adr_i[29]
port 335 nsew signal input
flabel metal3 s 200 13384 800 13608 0 FreeSans 896 0 0 0 wbs_adr_i[2]
port 336 nsew signal input
flabel metal3 s 200 46984 800 47208 0 FreeSans 896 0 0 0 wbs_adr_i[30]
port 337 nsew signal input
flabel metal3 s 119200 51016 119800 51240 0 FreeSans 896 0 0 0 wbs_adr_i[31]
port 338 nsew signal input
flabel metal2 s 93352 200 93576 800 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 339 nsew signal input
flabel metal2 s 92680 119200 92904 119800 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 340 nsew signal input
flabel metal2 s 89992 200 90216 800 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 341 nsew signal input
flabel metal3 s 200 57736 800 57960 0 FreeSans 896 0 0 0 wbs_adr_i[6]
port 342 nsew signal input
flabel metal2 s 5320 200 5544 800 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 343 nsew signal input
flabel metal3 s 119200 -56 119800 168 0 FreeSans 896 0 0 0 wbs_adr_i[8]
port 344 nsew signal input
flabel metal3 s 119200 32200 119800 32424 0 FreeSans 896 0 0 0 wbs_adr_i[9]
port 345 nsew signal input
flabel metal2 s 38248 119200 38472 119800 0 FreeSans 896 90 0 0 wbs_cyc_i
port 346 nsew signal input
flabel metal3 s 119200 104104 119800 104328 0 FreeSans 896 0 0 0 wbs_dat_i[0]
port 347 nsew signal input
flabel metal3 s 200 92680 800 92904 0 FreeSans 896 0 0 0 wbs_dat_i[10]
port 348 nsew signal input
flabel metal3 s 200 101416 800 101640 0 FreeSans 896 0 0 0 wbs_dat_i[11]
port 349 nsew signal input
flabel metal3 s 200 96712 800 96936 0 FreeSans 896 0 0 0 wbs_dat_i[12]
port 350 nsew signal input
flabel metal2 s 3976 200 4200 800 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 351 nsew signal input
flabel metal3 s 200 24808 800 25032 0 FreeSans 896 0 0 0 wbs_dat_i[14]
port 352 nsew signal input
flabel metal3 s 119200 62440 119800 62664 0 FreeSans 896 0 0 0 wbs_dat_i[15]
port 353 nsew signal input
flabel metal2 s 69160 200 69384 800 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 354 nsew signal input
flabel metal2 s 81928 119200 82152 119800 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 355 nsew signal input
flabel metal2 s 111496 119200 111720 119800 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 356 nsew signal input
flabel metal2 s 5992 119200 6216 119800 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 357 nsew signal input
flabel metal2 s 18088 200 18312 800 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 358 nsew signal input
flabel metal3 s 200 29512 800 29736 0 FreeSans 896 0 0 0 wbs_dat_i[20]
port 359 nsew signal input
flabel metal2 s 114856 119200 115080 119800 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 360 nsew signal input
flabel metal3 s 200 71176 800 71400 0 FreeSans 896 0 0 0 wbs_dat_i[22]
port 361 nsew signal input
flabel metal3 s 119200 94024 119800 94248 0 FreeSans 896 0 0 0 wbs_dat_i[23]
port 362 nsew signal input
flabel metal3 s 119200 39592 119800 39816 0 FreeSans 896 0 0 0 wbs_dat_i[24]
port 363 nsew signal input
flabel metal2 s 83272 200 83496 800 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 364 nsew signal input
flabel metal2 s 99400 119200 99624 119800 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 365 nsew signal input
flabel metal2 s 28840 119200 29064 119800 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 366 nsew signal input
flabel metal2 s 37576 200 37800 800 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 367 nsew signal input
flabel metal3 s 119200 73192 119800 73416 0 FreeSans 896 0 0 0 wbs_dat_i[29]
port 368 nsew signal input
flabel metal2 s 98056 200 98280 800 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 369 nsew signal input
flabel metal3 s 119200 35560 119800 35784 0 FreeSans 896 0 0 0 wbs_dat_i[30]
port 370 nsew signal input
flabel metal3 s 200 63112 800 63336 0 FreeSans 896 0 0 0 wbs_dat_i[31]
port 371 nsew signal input
flabel metal3 s 119200 4648 119800 4872 0 FreeSans 896 0 0 0 wbs_dat_i[3]
port 372 nsew signal input
flabel metal2 s 19432 200 19656 800 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 373 nsew signal input
flabel metal2 s 59752 200 59976 800 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 374 nsew signal input
flabel metal3 s 119200 52360 119800 52584 0 FreeSans 896 0 0 0 wbs_dat_i[6]
port 375 nsew signal input
flabel metal2 s 94696 119200 94920 119800 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 376 nsew signal input
flabel metal3 s 119200 107464 119800 107688 0 FreeSans 896 0 0 0 wbs_dat_i[8]
port 377 nsew signal input
flabel metal3 s 119200 5992 119800 6216 0 FreeSans 896 0 0 0 wbs_dat_i[9]
port 378 nsew signal input
flabel metal3 s 200 24136 800 24360 0 FreeSans 896 0 0 0 wbs_dat_o[0]
port 379 nsew signal tristate
flabel metal3 s 119200 68488 119800 68712 0 FreeSans 896 0 0 0 wbs_dat_o[10]
port 380 nsew signal tristate
flabel metal2 s 1960 200 2184 800 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 381 nsew signal tristate
flabel metal3 s 119200 110152 119800 110376 0 FreeSans 896 0 0 0 wbs_dat_o[12]
port 382 nsew signal tristate
flabel metal2 s 90664 119200 90888 119800 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 383 nsew signal tristate
flabel metal3 s 119200 14056 119800 14280 0 FreeSans 896 0 0 0 wbs_dat_o[14]
port 384 nsew signal tristate
flabel metal2 s 85960 119200 86184 119800 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 385 nsew signal tristate
flabel metal3 s 200 33544 800 33768 0 FreeSans 896 0 0 0 wbs_dat_o[16]
port 386 nsew signal tristate
flabel metal3 s 200 37576 800 37800 0 FreeSans 896 0 0 0 wbs_dat_o[17]
port 387 nsew signal tristate
flabel metal2 s 80584 200 80808 800 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 388 nsew signal tristate
flabel metal2 s -56 200 168 800 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 389 nsew signal tristate
flabel metal2 s 94696 200 94920 800 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 390 nsew signal tristate
flabel metal3 s 200 56392 800 56616 0 FreeSans 896 0 0 0 wbs_dat_o[20]
port 391 nsew signal tristate
flabel metal3 s 200 104104 800 104328 0 FreeSans 896 0 0 0 wbs_dat_o[21]
port 392 nsew signal tristate
flabel metal2 s 32200 119200 32424 119800 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 393 nsew signal tristate
flabel metal3 s 200 38920 800 39144 0 FreeSans 896 0 0 0 wbs_dat_o[23]
port 394 nsew signal tristate
flabel metal2 s 24808 200 25032 800 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 395 nsew signal tristate
flabel metal2 s 8680 200 8904 800 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 396 nsew signal tristate
flabel metal2 s 62440 119200 62664 119800 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 397 nsew signal tristate
flabel metal2 s 34888 119200 35112 119800 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 398 nsew signal tristate
flabel metal2 s 64456 200 64680 800 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 399 nsew signal tristate
flabel metal2 s 83272 119200 83496 119800 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 400 nsew signal tristate
flabel metal3 s 119200 33544 119800 33768 0 FreeSans 896 0 0 0 wbs_dat_o[2]
port 401 nsew signal tristate
flabel metal3 s 200 78568 800 78792 0 FreeSans 896 0 0 0 wbs_dat_o[30]
port 402 nsew signal tristate
flabel metal3 s 119200 92680 119800 92904 0 FreeSans 896 0 0 0 wbs_dat_o[31]
port 403 nsew signal tristate
flabel metal2 s 26152 200 26376 800 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 404 nsew signal tristate
flabel metal2 s 46312 200 46536 800 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 405 nsew signal tristate
flabel metal3 s 200 10024 800 10248 0 FreeSans 896 0 0 0 wbs_dat_o[5]
port 406 nsew signal tristate
flabel metal3 s 119200 89320 119800 89544 0 FreeSans 896 0 0 0 wbs_dat_o[6]
port 407 nsew signal tristate
flabel metal2 s 72520 200 72744 800 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 408 nsew signal tristate
flabel metal2 s 78568 119200 78792 119800 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 409 nsew signal tristate
flabel metal2 s 77896 119200 78120 119800 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 410 nsew signal tristate
flabel metal3 s 200 110824 800 111048 0 FreeSans 896 0 0 0 wbs_sel_i[0]
port 411 nsew signal input
flabel metal2 s 12712 119200 12936 119800 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 412 nsew signal input
flabel metal2 s 86632 200 86856 800 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 413 nsew signal input
flabel metal3 s 200 26152 800 26376 0 FreeSans 896 0 0 0 wbs_sel_i[3]
port 414 nsew signal input
flabel metal3 s 200 99400 800 99624 0 FreeSans 896 0 0 0 wbs_stb_i
port 415 nsew signal input
flabel metal3 s 119200 59080 119800 59304 0 FreeSans 896 0 0 0 wbs_we_i
port 416 nsew signal input
rlabel metal1 59976 116816 59976 116816 0 vdd
rlabel metal1 59976 116032 59976 116032 0 vss
rlabel metal3 47376 64568 47376 64568 0 _000_
rlabel metal2 47096 50064 47096 50064 0 _001_
rlabel metal2 92064 21672 92064 21672 0 _002_
rlabel metal2 115976 34440 115976 34440 0 _003_
rlabel metal3 45864 21672 45864 21672 0 _004_
rlabel metal3 46760 20888 46760 20888 0 _005_
rlabel metal2 46872 25032 46872 25032 0 _006_
rlabel metal2 115304 65632 115304 65632 0 _007_
rlabel metal2 70112 50008 70112 50008 0 _008_
rlabel metal2 78120 67816 78120 67816 0 _009_
rlabel metal2 75040 67144 75040 67144 0 _010_
rlabel metal2 66360 64904 66360 64904 0 _011_
rlabel metal2 46088 62440 46088 62440 0 _012_
rlabel metal2 117096 67396 117096 67396 0 _013_
rlabel metal2 72072 66976 72072 66976 0 _014_
rlabel metal2 71176 51800 71176 51800 0 _015_
rlabel metal2 69608 64904 69608 64904 0 _016_
rlabel metal3 46648 34216 46648 34216 0 _017_
rlabel metal2 53816 38780 53816 38780 0 _018_
rlabel metal2 78344 22568 78344 22568 0 _019_
rlabel metal2 46984 28168 46984 28168 0 _020_
rlabel metal3 46648 56168 46648 56168 0 _021_
rlabel metal3 46312 65576 46312 65576 0 _022_
rlabel metal2 47992 64232 47992 64232 0 _023_
rlabel metal3 47264 47544 47264 47544 0 _024_
rlabel metal2 47992 40712 47992 40712 0 _025_
rlabel metal2 47656 45976 47656 45976 0 _026_
rlabel metal2 61768 66528 61768 66528 0 _027_
rlabel metal3 49056 66360 49056 66360 0 _028_
rlabel metal2 61880 37688 61880 37688 0 _029_
rlabel metal3 72184 60984 72184 60984 0 _030_
rlabel metal2 50344 62776 50344 62776 0 _031_
rlabel metal2 72240 62552 72240 62552 0 _032_
rlabel metal2 61488 49112 61488 49112 0 _033_
rlabel metal3 55552 45976 55552 45976 0 _034_
rlabel metal2 64680 49224 64680 49224 0 _035_
rlabel metal2 59976 47152 59976 47152 0 _036_
rlabel metal3 58968 44408 58968 44408 0 _037_
rlabel metal2 61768 42448 61768 42448 0 _038_
rlabel metal2 64120 47096 64120 47096 0 _039_
rlabel metal3 66024 56952 66024 56952 0 _040_
rlabel metal2 65800 60312 65800 60312 0 _041_
rlabel metal3 61712 62328 61712 62328 0 _042_
rlabel metal2 63728 66360 63728 66360 0 _043_
rlabel metal2 54264 63504 54264 63504 0 _044_
rlabel metal2 53704 66696 53704 66696 0 _045_
rlabel metal2 58296 66640 58296 66640 0 _046_
rlabel metal2 52920 59920 52920 59920 0 _047_
rlabel metal3 59192 63896 59192 63896 0 _048_
rlabel metal3 60200 53928 60200 53928 0 _049_
rlabel metal2 55048 55272 55048 55272 0 _050_
rlabel metal2 64008 54040 64008 54040 0 _051_
rlabel metal3 49448 55496 49448 55496 0 _052_
rlabel metal3 53928 41272 53928 41272 0 _053_
rlabel metal3 54712 43624 54712 43624 0 _054_
rlabel metal2 51016 40656 51016 40656 0 _055_
rlabel metal2 68600 53648 68600 53648 0 _056_
rlabel metal2 68712 47432 68712 47432 0 _057_
rlabel metal2 51184 47544 51184 47544 0 _058_
rlabel metal3 49392 58520 49392 58520 0 _059_
rlabel metal3 48608 52360 48608 52360 0 _060_
rlabel metal2 50904 46256 50904 46256 0 _061_
rlabel metal2 70168 54040 70168 54040 0 _062_
rlabel metal3 70280 56952 70280 56952 0 _063_
rlabel metal2 67648 62216 67648 62216 0 _064_
rlabel metal2 63448 49672 63448 49672 0 _065_
rlabel metal2 62216 49112 62216 49112 0 _066_
rlabel metal3 40320 99176 40320 99176 0 _067_
rlabel metal2 43400 54040 43400 54040 0 _068_
rlabel metal3 68432 47320 68432 47320 0 _069_
rlabel metal2 48496 49112 48496 49112 0 _070_
rlabel metal2 59976 48888 59976 48888 0 _071_
rlabel metal2 60704 52360 60704 52360 0 _072_
rlabel metal2 47768 28952 47768 28952 0 _073_
rlabel metal3 47712 22456 47712 22456 0 _074_
rlabel metal3 46312 49784 46312 49784 0 _075_
rlabel metal3 48832 62440 48832 62440 0 _076_
rlabel metal3 47656 49896 47656 49896 0 _077_
rlabel metal2 91224 21616 91224 21616 0 _078_
rlabel metal2 116144 32760 116144 32760 0 _079_
rlabel metal2 44296 21840 44296 21840 0 _080_
rlabel metal2 45640 21644 45640 21644 0 _081_
rlabel metal2 46872 23800 46872 23800 0 _082_
rlabel metal2 45696 24136 45696 24136 0 _083_
rlabel metal3 114632 66248 114632 66248 0 _084_
rlabel metal3 68992 62888 68992 62888 0 _085_
rlabel metal3 71344 49672 71344 49672 0 _086_
rlabel metal2 77560 67508 77560 67508 0 _087_
rlabel metal2 74872 67144 74872 67144 0 _088_
rlabel metal2 66472 63784 66472 63784 0 _089_
rlabel metal2 66696 64176 66696 64176 0 _090_
rlabel metal2 45752 61152 45752 61152 0 _091_
rlabel metal2 117488 67816 117488 67816 0 _092_
rlabel metal2 71400 67480 71400 67480 0 _093_
rlabel metal2 71176 51296 71176 51296 0 _094_
rlabel metal3 71848 51352 71848 51352 0 _095_
rlabel metal2 67648 64568 67648 64568 0 _096_
rlabel metal3 70280 64568 70280 64568 0 _097_
rlabel metal2 46032 33544 46032 33544 0 _098_
rlabel metal3 53928 37464 53928 37464 0 _099_
rlabel metal3 78120 23128 78120 23128 0 _100_
rlabel metal2 45752 27888 45752 27888 0 _101_
rlabel metal2 46424 56168 46424 56168 0 _102_
rlabel metal2 45640 65576 45640 65576 0 _103_
rlabel metal2 48216 64512 48216 64512 0 _104_
rlabel metal3 49000 63784 49000 63784 0 _105_
rlabel metal2 47096 48552 47096 48552 0 _106_
rlabel metal2 47320 48160 47320 48160 0 _107_
rlabel metal2 48104 40488 48104 40488 0 _108_
rlabel metal3 48776 46648 48776 46648 0 _109_
rlabel metal2 47824 45304 47824 45304 0 _110_
rlabel metal2 61544 66920 61544 66920 0 _111_
rlabel metal3 49056 67032 49056 67032 0 _112_
rlabel metal2 61712 38584 61712 38584 0 _113_
rlabel metal2 70280 61152 70280 61152 0 _114_
rlabel metal3 72968 60648 72968 60648 0 _115_
rlabel metal2 69440 61544 69440 61544 0 _116_
rlabel metal2 50568 62440 50568 62440 0 _117_
rlabel metal2 70952 61488 70952 61488 0 _118_
rlabel metal3 72968 62328 72968 62328 0 _119_
rlabel metal2 56392 51744 56392 51744 0 _120_
rlabel via2 65016 50568 65016 50568 0 _121_
rlabel metal2 67032 48048 67032 48048 0 _122_
rlabel metal2 63112 47768 63112 47768 0 _123_
rlabel metal2 65800 48440 65800 48440 0 _124_
rlabel metal2 56728 52808 56728 52808 0 _125_
rlabel metal2 62216 58688 62216 58688 0 _126_
rlabel metal2 63112 52416 63112 52416 0 _127_
rlabel metal2 56112 48888 56112 48888 0 _128_
rlabel metal2 56448 52360 56448 52360 0 _129_
rlabel metal2 62888 59696 62888 59696 0 _130_
rlabel metal2 55888 60536 55888 60536 0 _131_
rlabel metal3 54432 62216 54432 62216 0 _132_
rlabel metal2 41720 55272 41720 55272 0 _133_
rlabel metal3 45024 55272 45024 55272 0 _134_
rlabel metal2 68432 56056 68432 56056 0 _135_
rlabel metal3 53368 55384 53368 55384 0 _136_
rlabel metal2 55048 54600 55048 54600 0 _137_
rlabel metal2 56280 53200 56280 53200 0 _138_
rlabel metal2 57904 65576 57904 65576 0 _139_
rlabel metal3 63560 65352 63560 65352 0 _140_
rlabel metal3 58856 60760 58856 60760 0 _141_
rlabel metal2 53816 64792 53816 64792 0 _142_
rlabel metal2 59752 57008 59752 57008 0 _143_
rlabel metal2 64008 43120 64008 43120 0 _144_
rlabel metal2 68040 44408 68040 44408 0 _145_
rlabel metal2 48888 43232 48888 43232 0 _146_
rlabel metal2 59192 42392 59192 42392 0 _147_
rlabel metal2 59864 43736 59864 43736 0 _148_
rlabel metal2 58968 55496 58968 55496 0 _149_
rlabel metal2 43344 52024 43344 52024 0 _150_
rlabel metal2 63672 55664 63672 55664 0 _151_
rlabel metal3 56392 45864 56392 45864 0 _152_
rlabel metal2 59192 55048 59192 55048 0 _153_
rlabel metal2 59696 58632 59696 58632 0 _154_
rlabel metal3 59024 58632 59024 58632 0 _155_
rlabel metal3 58744 58408 58744 58408 0 _156_
rlabel metal2 58968 58744 58968 58744 0 _157_
rlabel metal2 59080 57176 59080 57176 0 _158_
rlabel metal2 56056 54376 56056 54376 0 _159_
rlabel metal2 56504 46872 56504 46872 0 _160_
rlabel metal3 65296 48888 65296 48888 0 _161_
rlabel metal2 61376 48888 61376 48888 0 _162_
rlabel metal2 64008 50960 64008 50960 0 _163_
rlabel metal3 65016 45192 65016 45192 0 _164_
rlabel metal2 55664 47432 55664 47432 0 _165_
rlabel metal2 56056 48216 56056 48216 0 _166_
rlabel metal2 56056 46984 56056 46984 0 _167_
rlabel metal3 63672 48216 63672 48216 0 _168_
rlabel metal2 63224 48496 63224 48496 0 _169_
rlabel metal3 63504 49112 63504 49112 0 _170_
rlabel metal2 64456 50344 64456 50344 0 _171_
rlabel metal3 60928 48104 60928 48104 0 _172_
rlabel metal2 59416 48216 59416 48216 0 _173_
rlabel metal2 58408 47656 58408 47656 0 _174_
rlabel metal3 59192 47656 59192 47656 0 _175_
rlabel metal3 58184 59976 58184 59976 0 _176_
rlabel metal3 57848 45080 57848 45080 0 _177_
rlabel metal3 59304 45080 59304 45080 0 _178_
rlabel metal2 58184 42728 58184 42728 0 _179_
rlabel metal3 64736 46760 64736 46760 0 _180_
rlabel metal2 58072 42392 58072 42392 0 _181_
rlabel metal2 59304 43456 59304 43456 0 _182_
rlabel metal2 59528 42168 59528 42168 0 _183_
rlabel metal3 60424 42616 60424 42616 0 _184_
rlabel metal2 64120 46256 64120 46256 0 _185_
rlabel metal2 62776 44744 62776 44744 0 _186_
rlabel metal2 63000 45416 63000 45416 0 _187_
rlabel metal3 63392 46648 63392 46648 0 _188_
rlabel metal2 63672 58072 63672 58072 0 _189_
rlabel metal2 69048 63672 69048 63672 0 _190_
rlabel metal2 64456 57008 64456 57008 0 _191_
rlabel metal3 64456 57064 64456 57064 0 _192_
rlabel metal3 64512 65576 64512 65576 0 _193_
rlabel metal2 56392 58968 56392 58968 0 _194_
rlabel metal2 57064 59696 57064 59696 0 _195_
rlabel metal2 62552 65352 62552 65352 0 _196_
rlabel metal3 64680 62328 64680 62328 0 _197_
rlabel metal2 63336 59584 63336 59584 0 _198_
rlabel metal2 56616 66360 56616 66360 0 _199_
rlabel metal2 63672 59976 63672 59976 0 _200_
rlabel metal2 63784 62720 63784 62720 0 _201_
rlabel metal3 64792 63896 64792 63896 0 _202_
rlabel metal2 63672 64232 63672 64232 0 _203_
rlabel metal2 62328 63000 62328 63000 0 _204_
rlabel metal2 61936 62888 61936 62888 0 _205_
rlabel metal3 60424 60760 60424 60760 0 _206_
rlabel metal2 63448 64904 63448 64904 0 _207_
rlabel metal2 63336 66696 63336 66696 0 _208_
rlabel metal2 63896 63504 63896 63504 0 _209_
rlabel metal2 55160 63112 55160 63112 0 _210_
rlabel metal2 55272 63112 55272 63112 0 _211_
rlabel metal3 55608 67144 55608 67144 0 _212_
rlabel metal2 55272 66528 55272 66528 0 _213_
rlabel metal3 54712 66136 54712 66136 0 _214_
rlabel metal2 56616 67592 56616 67592 0 _215_
rlabel metal2 57064 67144 57064 67144 0 _216_
rlabel metal2 57960 66024 57960 66024 0 _217_
rlabel metal2 62888 58352 62888 58352 0 _218_
rlabel metal2 57624 62188 57624 62188 0 _219_
rlabel metal2 56056 59248 56056 59248 0 _220_
rlabel metal2 53928 61824 53928 61824 0 _221_
rlabel metal2 55384 60256 55384 60256 0 _222_
rlabel metal2 54376 60144 54376 60144 0 _223_
rlabel metal2 58520 62720 58520 62720 0 _224_
rlabel metal2 58184 63280 58184 63280 0 _225_
rlabel metal3 58520 52808 58520 52808 0 _226_
rlabel metal3 59528 48888 59528 48888 0 _227_
rlabel metal2 57736 51408 57736 51408 0 _228_
rlabel metal3 49056 42728 49056 42728 0 _229_
rlabel metal2 56504 55272 56504 55272 0 _230_
rlabel metal2 58072 53760 58072 53760 0 _231_
rlabel metal2 66472 44912 66472 44912 0 _232_
rlabel metal2 57960 53480 57960 53480 0 _233_
rlabel metal2 53032 54768 53032 54768 0 _234_
rlabel metal3 55048 55944 55048 55944 0 _235_
rlabel metal2 57624 57288 57624 57288 0 _236_
rlabel metal2 60200 56896 60200 56896 0 _237_
rlabel metal3 54376 56056 54376 56056 0 _238_
rlabel metal2 55048 55888 55048 55888 0 _239_
rlabel metal2 61768 55608 61768 55608 0 _240_
rlabel metal3 63000 55048 63000 55048 0 _241_
rlabel metal3 48104 50232 48104 50232 0 _242_
rlabel metal2 48440 54264 48440 54264 0 _243_
rlabel metal2 51800 54544 51800 54544 0 _244_
rlabel metal2 50120 55664 50120 55664 0 _245_
rlabel metal2 50008 55888 50008 55888 0 _246_
rlabel metal2 52136 43064 52136 43064 0 _247_
rlabel metal2 53088 42504 53088 42504 0 _248_
rlabel metal3 52976 44072 52976 44072 0 _249_
rlabel metal2 52920 51688 52920 51688 0 _250_
rlabel metal2 49560 43848 49560 43848 0 _251_
rlabel metal2 54264 44632 54264 44632 0 _252_
rlabel metal2 67144 44016 67144 44016 0 _253_
rlabel metal2 50232 43064 50232 43064 0 _254_
rlabel metal2 50680 40432 50680 40432 0 _255_
rlabel metal2 67368 56448 67368 56448 0 _256_
rlabel metal2 48944 48440 48944 48440 0 _257_
rlabel metal2 67200 52248 67200 52248 0 _258_
rlabel metal2 67928 55440 67928 55440 0 _259_
rlabel metal2 54544 50008 54544 50008 0 _260_
rlabel metal2 54264 50736 54264 50736 0 _261_
rlabel metal3 49896 49000 49896 49000 0 _262_
rlabel metal2 66920 50008 66920 50008 0 _263_
rlabel metal2 67256 48944 67256 48944 0 _264_
rlabel metal2 49504 49000 49504 49000 0 _265_
rlabel metal3 67816 48328 67816 48328 0 _266_
rlabel metal2 50456 50736 50456 50736 0 _267_
rlabel metal2 51576 50232 51576 50232 0 _268_
rlabel metal2 50344 50848 50344 50848 0 _269_
rlabel metal3 51464 48328 51464 48328 0 _270_
rlabel metal2 50232 48944 50232 48944 0 _271_
rlabel metal2 50456 50204 50456 50204 0 _272_
rlabel metal2 50960 50344 50960 50344 0 _273_
rlabel metal2 49784 60312 49784 60312 0 _274_
rlabel metal2 49560 59528 49560 59528 0 _275_
rlabel metal2 49784 53760 49784 53760 0 _276_
rlabel metal2 50064 52360 50064 52360 0 _277_
rlabel metal2 50232 52976 50232 52976 0 _278_
rlabel metal2 68824 50960 68824 50960 0 _279_
rlabel metal3 48272 53928 48272 53928 0 _280_
rlabel metal2 49560 52920 49560 52920 0 _281_
rlabel metal2 52136 49392 52136 49392 0 _282_
rlabel metal2 50008 49280 50008 49280 0 _283_
rlabel metal2 50344 47432 50344 47432 0 _284_
rlabel metal2 70336 57624 70336 57624 0 _285_
rlabel metal2 70000 55272 70000 55272 0 _286_
rlabel metal2 70392 54488 70392 54488 0 _287_
rlabel metal2 70896 57848 70896 57848 0 _288_
rlabel metal2 69608 60872 69608 60872 0 _289_
rlabel metal2 70728 59864 70728 59864 0 _290_
rlabel metal2 69496 58016 69496 58016 0 _291_
rlabel metal2 69720 56952 69720 56952 0 _292_
rlabel metal2 68376 59584 68376 59584 0 _293_
rlabel metal2 68712 60200 68712 60200 0 _294_
rlabel metal2 67928 60200 67928 60200 0 _295_
rlabel metal2 66304 59080 66304 59080 0 _296_
rlabel metal2 67536 60872 67536 60872 0 _297_
rlabel metal2 69384 28336 69384 28336 0 clknet_0_wb_clk_i
rlabel metal2 47768 27776 47768 27776 0 clknet_3_0__leaf_wb_clk_i
rlabel metal3 69944 30072 69944 30072 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 49896 41496 49896 41496 0 clknet_3_2__leaf_wb_clk_i
rlabel metal3 63392 45752 63392 45752 0 clknet_3_3__leaf_wb_clk_i
rlabel metal3 48552 65464 48552 65464 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 67872 49112 67872 49112 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 50232 66304 50232 66304 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 74984 62104 74984 62104 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 3528 117530 3528 117530 0 io_oeb[0]
rlabel metal3 1358 82152 1358 82152 0 io_oeb[10]
rlabel metal3 1358 75432 1358 75432 0 io_oeb[11]
rlabel metal3 1358 90216 1358 90216 0 io_oeb[12]
rlabel metal2 102984 2198 102984 2198 0 io_oeb[13]
rlabel metal2 117656 2478 117656 2478 0 io_oeb[14]
rlabel metal2 65240 116760 65240 116760 0 io_oeb[15]
rlabel metal3 1358 69272 1358 69272 0 io_oeb[16]
rlabel metal2 11760 115528 11760 115528 0 io_oeb[17]
rlabel metal3 1358 94920 1358 94920 0 io_oeb[18]
rlabel metal2 48552 2198 48552 2198 0 io_oeb[19]
rlabel metal2 115528 9744 115528 9744 0 io_oeb[1]
rlabel metal2 102424 2464 102424 2464 0 io_oeb[20]
rlabel metal2 11480 2198 11480 2198 0 io_oeb[21]
rlabel metal2 115528 30632 115528 30632 0 io_oeb[22]
rlabel metal3 1358 11592 1358 11592 0 io_oeb[23]
rlabel metal2 115528 27104 115528 27104 0 io_oeb[24]
rlabel metal2 42280 2478 42280 2478 0 io_oeb[25]
rlabel metal2 99624 798 99624 798 0 io_oeb[26]
rlabel metal3 1358 80136 1358 80136 0 io_oeb[27]
rlabel metal3 1358 112392 1358 112392 0 io_oeb[28]
rlabel metal3 25200 116536 25200 116536 0 io_oeb[29]
rlabel metal2 77448 798 77448 798 0 io_oeb[2]
rlabel metal3 1302 4200 1302 4200 0 io_oeb[30]
rlabel metal2 115416 83552 115416 83552 0 io_oeb[31]
rlabel metal2 115528 19152 115528 19152 0 io_oeb[32]
rlabel metal3 1358 98280 1358 98280 0 io_oeb[33]
rlabel metal3 1358 46536 1358 46536 0 io_oeb[34]
rlabel metal3 68264 116536 68264 116536 0 io_oeb[35]
rlabel metal2 112392 2142 112392 2142 0 io_oeb[36]
rlabel metal2 115528 40880 115528 40880 0 io_oeb[3]
rlabel metal2 168 118594 168 118594 0 io_oeb[4]
rlabel metal3 117418 115528 117418 115528 0 io_oeb[5]
rlabel metal2 58296 116480 58296 116480 0 io_oeb[6]
rlabel metal2 115528 7112 115528 7112 0 io_oeb[7]
rlabel metal2 115528 48832 115528 48832 0 io_oeb[8]
rlabel metal2 115528 47992 115528 47992 0 io_oeb[9]
rlabel metal3 1358 23016 1358 23016 0 io_out[0]
rlabel metal2 115864 115136 115864 115136 0 io_out[10]
rlabel metal3 117586 105672 117586 105672 0 io_out[11]
rlabel metal2 117880 116984 117880 116984 0 io_out[12]
rlabel metal3 1358 88872 1358 88872 0 io_out[13]
rlabel metal2 47208 2478 47208 2478 0 io_out[14]
rlabel metal3 117586 99624 117586 99624 0 io_out[15]
rlabel metal2 13608 2478 13608 2478 0 io_out[16]
rlabel metal2 100968 2086 100968 2086 0 io_out[17]
rlabel metal2 78792 2478 78792 2478 0 io_out[18]
rlabel metal2 8008 2198 8008 2198 0 io_out[19]
rlabel metal2 82152 2478 82152 2478 0 io_out[1]
rlabel metal2 54600 2478 54600 2478 0 io_out[20]
rlabel metal2 40488 2870 40488 2870 0 io_out[21]
rlabel metal3 1358 16296 1358 16296 0 io_out[22]
rlabel metal3 88648 116536 88648 116536 0 io_out[23]
rlabel metal2 55720 117418 55720 117418 0 io_out[24]
rlabel metal2 50456 2086 50456 2086 0 io_out[25]
rlabel metal2 86632 116760 86632 116760 0 io_out[26]
rlabel metal2 88872 2086 88872 2086 0 io_out[27]
rlabel metal2 77560 115640 77560 115640 0 io_out[28]
rlabel metal2 113736 3262 113736 3262 0 io_out[29]
rlabel metal2 110376 117530 110376 117530 0 io_out[2]
rlabel metal3 117586 25704 117586 25704 0 io_out[30]
rlabel metal3 101360 115528 101360 115528 0 io_out[31]
rlabel metal3 117586 86184 117586 86184 0 io_out[3]
rlabel metal3 2254 3528 2254 3528 0 io_out[4]
rlabel metal3 1358 5544 1358 5544 0 io_out[5]
rlabel metal3 1358 68040 1358 68040 0 io_out[6]
rlabel metal3 76216 116536 76216 116536 0 io_out[7]
rlabel metal2 31080 798 31080 798 0 io_out[8]
rlabel metal3 1358 61320 1358 61320 0 io_out[9]
rlabel metal3 60256 116536 60256 116536 0 la_data_in[32]
rlabel metal3 118202 102088 118202 102088 0 la_data_in[33]
rlabel metal2 37016 117922 37016 117922 0 la_data_in[34]
rlabel metal2 49616 116536 49616 116536 0 la_data_in[35]
rlabel metal2 116984 64960 116984 64960 0 la_data_in[36]
rlabel metal2 41552 3416 41552 3416 0 la_data_in[37]
rlabel metal2 57680 3416 57680 3416 0 la_data_in[38]
rlabel metal3 1246 40488 1246 40488 0 la_data_in[39]
rlabel metal2 114520 2464 114520 2464 0 la_data_in[40]
rlabel metal2 1848 113456 1848 113456 0 la_data_in[41]
rlabel metal2 116872 87136 116872 87136 0 la_data_in[42]
rlabel metal3 74592 3416 74592 3416 0 la_data_in[43]
rlabel metal2 56224 116536 56224 116536 0 la_data_in[44]
rlabel metal2 15736 116872 15736 116872 0 la_data_in[45]
rlabel metal2 10024 116536 10024 116536 0 la_data_in[46]
rlabel metal3 47320 116312 47320 116312 0 la_data_in[47]
rlabel metal2 55272 2086 55272 2086 0 la_data_in[48]
rlabel metal3 1302 62552 1302 62552 0 la_data_in[49]
rlabel metal2 1960 37240 1960 37240 0 la_data_in[50]
rlabel metal2 1848 31892 1848 31892 0 la_data_in[51]
rlabel metal3 1470 35784 1470 35784 0 la_data_in[52]
rlabel metal2 117880 3864 117880 3864 0 la_data_in[53]
rlabel metal2 44072 3808 44072 3808 0 la_data_in[54]
rlabel metal3 116872 109144 116872 109144 0 la_data_in[55]
rlabel metal3 21280 3416 21280 3416 0 la_data_in[56]
rlabel metal2 31472 116312 31472 116312 0 la_data_in[57]
rlabel metal2 45080 117922 45080 117922 0 la_data_in[58]
rlabel metal2 70504 4200 70504 4200 0 la_data_in[59]
rlabel metal2 24696 2072 24696 2072 0 la_data_in[60]
rlabel metal2 116872 43288 116872 43288 0 la_data_in[61]
rlabel metal2 35392 116312 35392 116312 0 la_data_in[62]
rlabel metal2 108752 115864 108752 115864 0 la_data_in[63]
rlabel metal2 33992 116032 33992 116032 0 la_data_out[0]
rlabel metal2 115528 50288 115528 50288 0 la_data_out[10]
rlabel metal3 1358 102984 1358 102984 0 la_data_out[11]
rlabel metal3 117418 66024 117418 66024 0 la_data_out[12]
rlabel metal2 60088 115696 60088 115696 0 la_data_out[13]
rlabel metal3 53648 116536 53648 116536 0 la_data_out[14]
rlabel metal2 63336 2086 63336 2086 0 la_data_out[15]
rlabel metal3 117586 55944 117586 55944 0 la_data_out[16]
rlabel metal3 116928 115192 116928 115192 0 la_data_out[17]
rlabel metal2 2072 116928 2072 116928 0 la_data_out[18]
rlabel metal3 117698 75432 117698 75432 0 la_data_out[19]
rlabel metal2 35560 2198 35560 2198 0 la_data_out[1]
rlabel metal3 117586 35112 117586 35112 0 la_data_out[20]
rlabel metal3 1358 21000 1358 21000 0 la_data_out[21]
rlabel metal3 117586 14952 117586 14952 0 la_data_out[22]
rlabel metal2 74200 115696 74200 115696 0 la_data_out[23]
rlabel metal3 117586 94920 117586 94920 0 la_data_out[24]
rlabel metal2 51912 2478 51912 2478 0 la_data_out[25]
rlabel metal3 1358 93576 1358 93576 0 la_data_out[26]
rlabel metal3 117586 54600 117586 54600 0 la_data_out[27]
rlabel metal3 1358 45192 1358 45192 0 la_data_out[28]
rlabel metal2 70616 117922 70616 117922 0 la_data_out[29]
rlabel metal2 115528 22400 115528 22400 0 la_data_out[2]
rlabel metal2 58408 2478 58408 2478 0 la_data_out[30]
rlabel metal3 65912 116536 65912 116536 0 la_data_out[31]
rlabel metal2 6888 798 6888 798 0 la_data_out[3]
rlabel metal3 2142 2184 2142 2184 0 la_data_out[4]
rlabel metal3 117586 8232 117586 8232 0 la_data_out[5]
rlabel metal2 115528 45584 115528 45584 0 la_data_out[6]
rlabel metal3 117586 84840 117586 84840 0 la_data_out[7]
rlabel metal3 117474 67368 117474 67368 0 la_data_out[8]
rlabel metal2 47992 115640 47992 115640 0 la_data_out[9]
rlabel metal3 1400 4424 1400 4424 0 la_oenb[32]
rlabel metal2 1960 116704 1960 116704 0 la_oenb[33]
rlabel metal2 62776 4256 62776 4256 0 la_oenb[34]
rlabel metal2 1848 51632 1848 51632 0 la_oenb[35]
rlabel metal2 1848 65744 1848 65744 0 la_oenb[36]
rlabel metal2 1960 34608 1960 34608 0 la_oenb[37]
rlabel metal2 43736 117530 43736 117530 0 la_oenb[38]
rlabel metal2 1960 76328 1960 76328 0 la_oenb[39]
rlabel metal2 53144 2086 53144 2086 0 la_oenb[40]
rlabel metal3 1358 59864 1358 59864 0 la_oenb[41]
rlabel metal2 95984 3416 95984 3416 0 la_oenb[42]
rlabel metal2 45304 3416 45304 3416 0 la_oenb[43]
rlabel metal3 1358 88088 1358 88088 0 la_oenb[44]
rlabel metal2 117096 58072 117096 58072 0 la_oenb[45]
rlabel metal2 117992 79856 117992 79856 0 la_oenb[46]
rlabel metal2 92624 4200 92624 4200 0 la_oenb[47]
rlabel metal2 41160 116704 41160 116704 0 la_oenb[48]
rlabel metal2 117320 5152 117320 5152 0 la_oenb[49]
rlabel metal2 81200 116536 81200 116536 0 la_oenb[50]
rlabel metal3 118202 61320 118202 61320 0 la_oenb[51]
rlabel metal2 91336 2086 91336 2086 0 la_oenb[52]
rlabel metal2 106904 117922 106904 117922 0 la_oenb[53]
rlabel metal2 116872 11928 116872 11928 0 la_oenb[54]
rlabel metal2 72128 114968 72128 114968 0 la_oenb[55]
rlabel metal2 110936 2086 110936 2086 0 la_oenb[56]
rlabel metal3 1302 58520 1302 58520 0 la_oenb[57]
rlabel metal2 14672 3416 14672 3416 0 la_oenb[58]
rlabel metal3 118090 60648 118090 60648 0 la_oenb[59]
rlabel metal2 117992 78400 117992 78400 0 la_oenb[60]
rlabel metal2 29456 3416 29456 3416 0 la_oenb[61]
rlabel metal3 115416 3416 115416 3416 0 la_oenb[62]
rlabel metal2 1848 21560 1848 21560 0 la_oenb[63]
rlabel metal2 61040 116536 61040 116536 0 net1
rlabel metal2 3360 113960 3360 113960 0 net10
rlabel metal2 14280 90104 14280 90104 0 net100
rlabel metal3 83384 24920 83384 24920 0 net101
rlabel metal2 3304 27216 3304 27216 0 net102
rlabel metal2 37912 99568 37912 99568 0 net103
rlabel metal2 114968 59584 114968 59584 0 net104
rlabel metal2 3976 115192 3976 115192 0 net105
rlabel metal2 2520 82264 2520 82264 0 net106
rlabel metal2 2520 75376 2520 75376 0 net107
rlabel metal2 2520 90104 2520 90104 0 net108
rlabel metal2 103880 3976 103880 3976 0 net109
rlabel metal2 74760 76608 74760 76608 0 net11
rlabel metal2 117096 4368 117096 4368 0 net110
rlabel metal2 63896 115584 63896 115584 0 net111
rlabel metal2 2520 69832 2520 69832 0 net112
rlabel metal2 10696 115696 10696 115696 0 net113
rlabel metal2 2632 94360 2632 94360 0 net114
rlabel metal2 48832 4872 48832 4872 0 net115
rlabel metal2 117096 9744 117096 9744 0 net116
rlabel metal2 101192 4368 101192 4368 0 net117
rlabel metal2 11536 4424 11536 4424 0 net118
rlabel metal2 117096 30240 117096 30240 0 net119
rlabel metal2 74200 32424 74200 32424 0 net12
rlabel metal2 2856 11704 2856 11704 0 net120
rlabel metal3 116648 26936 116648 26936 0 net121
rlabel metal2 42728 4592 42728 4592 0 net122
rlabel metal2 99512 4200 99512 4200 0 net123
rlabel metal2 2520 80080 2520 80080 0 net124
rlabel metal2 2520 112784 2520 112784 0 net125
rlabel metal2 23576 116144 23576 116144 0 net126
rlabel metal2 77336 3976 77336 3976 0 net127
rlabel metal2 2520 4200 2520 4200 0 net128
rlabel metal3 116648 83384 116648 83384 0 net129
rlabel metal3 58856 116536 58856 116536 0 net13
rlabel metal2 117096 19152 117096 19152 0 net130
rlabel metal2 2856 98672 2856 98672 0 net131
rlabel metal2 2856 46928 2856 46928 0 net132
rlabel metal2 67256 116424 67256 116424 0 net133
rlabel metal3 112728 4872 112728 4872 0 net134
rlabel metal2 117096 40880 117096 40880 0 net135
rlabel metal2 3080 115920 3080 115920 0 net136
rlabel metal2 117096 114912 117096 114912 0 net137
rlabel metal2 57848 115192 57848 115192 0 net138
rlabel metal2 117096 7056 117096 7056 0 net139
rlabel metal2 16800 116536 16800 116536 0 net14
rlabel metal2 117096 48720 117096 48720 0 net140
rlabel metal2 117096 47768 117096 47768 0 net141
rlabel metal2 3080 23072 3080 23072 0 net142
rlabel metal2 117320 50288 117320 50288 0 net143
rlabel metal2 45920 62216 45920 62216 0 net144
rlabel metal2 117320 67480 117320 67480 0 net145
rlabel metal3 4312 88984 4312 88984 0 net146
rlabel metal3 49504 5208 49504 5208 0 net147
rlabel metal2 114744 99960 114744 99960 0 net148
rlabel metal3 48160 33432 48160 33432 0 net149
rlabel metal2 21000 89936 21000 89936 0 net15
rlabel metal2 100296 3864 100296 3864 0 net150
rlabel metal3 78624 4312 78624 4312 0 net151
rlabel metal2 47376 27160 47376 27160 0 net152
rlabel metal3 54432 4984 54432 4984 0 net153
rlabel metal3 57008 4312 57008 4312 0 net154
rlabel metal2 47264 64456 47264 64456 0 net155
rlabel metal3 3304 16856 3304 16856 0 net156
rlabel metal3 72072 115640 72072 115640 0 net157
rlabel metal3 71568 94360 71568 94360 0 net158
rlabel metal2 50680 4480 50680 4480 0 net159
rlabel metal2 48104 116368 48104 116368 0 net16
rlabel metal2 48664 93632 48664 93632 0 net160
rlabel metal2 49560 67816 49560 67816 0 net161
rlabel metal2 76888 115584 76888 115584 0 net162
rlabel metal3 70840 63896 70840 63896 0 net163
rlabel metal2 116648 24696 116648 24696 0 net164
rlabel metal2 68432 4536 68432 4536 0 net165
rlabel metal2 70168 115472 70168 115472 0 net166
rlabel metal2 46312 4480 46312 4480 0 net167
rlabel metal2 5656 4816 5656 4816 0 net168
rlabel metal3 3304 5880 3304 5880 0 net169
rlabel metal2 54824 3640 54824 3640 0 net17
rlabel metal2 3640 68432 3640 68432 0 net170
rlabel metal2 76272 116424 76272 116424 0 net171
rlabel metal2 78232 66192 78232 66192 0 net172
rlabel metal2 46088 68544 46088 68544 0 net173
rlabel metal2 34888 114744 34888 114744 0 net174
rlabel metal2 117096 50512 117096 50512 0 net175
rlabel metal2 3080 103040 3080 103040 0 net176
rlabel metal2 116200 67508 116200 67508 0 net177
rlabel metal2 59192 115304 59192 115304 0 net178
rlabel metal2 52752 116200 52752 116200 0 net179
rlabel metal2 3416 63224 3416 63224 0 net18
rlabel metal2 74088 41636 74088 41636 0 net180
rlabel metal2 114968 56112 114968 56112 0 net181
rlabel metal2 117432 67592 117432 67592 0 net182
rlabel metal3 3416 114856 3416 114856 0 net183
rlabel metal3 114688 75656 114688 75656 0 net184
rlabel metal2 54488 4480 54488 4480 0 net185
rlabel metal2 95704 35168 95704 35168 0 net186
rlabel metal2 3640 21392 3640 21392 0 net187
rlabel metal2 114968 15344 114968 15344 0 net188
rlabel metal2 72632 115696 72632 115696 0 net189
rlabel metal2 3360 37128 3360 37128 0 net19
rlabel metal2 114520 94696 114520 94696 0 net190
rlabel metal2 51016 4368 51016 4368 0 net191
rlabel metal2 3080 93632 3080 93632 0 net192
rlabel metal2 114408 54824 114408 54824 0 net193
rlabel metal2 3080 45752 3080 45752 0 net194
rlabel metal2 71232 115528 71232 115528 0 net195
rlabel metal2 116648 22344 116648 22344 0 net196
rlabel metal2 59528 4368 59528 4368 0 net197
rlabel metal2 68712 115976 68712 115976 0 net198
rlabel metal2 8232 4256 8232 4256 0 net199
rlabel metal3 85904 102424 85904 102424 0 net2
rlabel metal3 19768 32424 19768 32424 0 net20
rlabel metal2 5992 3976 5992 3976 0 net200
rlabel metal3 114744 8232 114744 8232 0 net201
rlabel metal2 117096 45584 117096 45584 0 net202
rlabel metal2 114744 85064 114744 85064 0 net203
rlabel metal2 114184 67928 114184 67928 0 net204
rlabel metal2 46984 115304 46984 115304 0 net205
rlabel metal2 91560 44744 91560 44744 0 net206
rlabel metal2 3080 24640 3080 24640 0 net207
rlabel metal3 114688 69384 114688 69384 0 net208
rlabel metal2 4984 4760 4984 4760 0 net209
rlabel metal2 37576 39144 37576 39144 0 net21
rlabel metal2 116424 68768 116424 68768 0 net210
rlabel metal2 92008 116312 92008 116312 0 net211
rlabel metal2 100296 32704 100296 32704 0 net212
rlabel metal2 72408 67676 72408 67676 0 net213
rlabel metal2 3080 34048 3080 34048 0 net214
rlabel metal2 3080 37912 3080 37912 0 net215
rlabel metal2 80752 3528 80752 3528 0 net216
rlabel metal2 3080 6552 3080 6552 0 net217
rlabel metal2 94808 3976 94808 3976 0 net218
rlabel metal2 3080 56728 3080 56728 0 net219
rlabel metal2 114968 4312 114968 4312 0 net22
rlabel metal2 3080 104608 3080 104608 0 net220
rlabel metal2 45864 63896 45864 63896 0 net221
rlabel metal2 3640 40432 3640 40432 0 net222
rlabel metal3 26656 5096 26656 5096 0 net223
rlabel metal2 10640 3528 10640 3528 0 net224
rlabel metal2 64176 67928 64176 67928 0 net225
rlabel metal2 49672 67396 49672 67396 0 net226
rlabel metal2 65184 3528 65184 3528 0 net227
rlabel metal2 74312 61320 74312 61320 0 net228
rlabel metal2 117208 33320 117208 33320 0 net229
rlabel metal2 45360 6328 45360 6328 0 net23
rlabel metal3 4704 78568 4704 78568 0 net230
rlabel metal3 114688 92904 114688 92904 0 net231
rlabel metal2 28168 4872 28168 4872 0 net232
rlabel metal2 46424 5208 46424 5208 0 net233
rlabel metal3 45696 23800 45696 23800 0 net234
rlabel metal2 116200 73080 116200 73080 0 net235
rlabel metal2 73304 4312 73304 4312 0 net236
rlabel metal2 78904 66248 78904 66248 0 net237
rlabel metal3 77504 68824 77504 68824 0 net238
rlabel metal3 3080 74984 3080 74984 0 net239
rlabel metal2 93240 82544 93240 82544 0 net24
rlabel metal2 2856 3920 2856 3920 0 net240
rlabel metal2 101416 4704 101416 4704 0 net241
rlabel metal2 76776 4536 76776 4536 0 net242
rlabel metal3 116480 114296 116480 114296 0 net243
rlabel metal3 1302 100968 1302 100968 0 net244
rlabel metal2 118104 38808 118104 38808 0 net245
rlabel metal2 80136 2030 80136 2030 0 net246
rlabel metal2 118104 78344 118104 78344 0 net247
rlabel metal2 28672 3304 28672 3304 0 net248
rlabel metal3 118104 112504 118104 112504 0 net249
rlabel metal2 22680 21728 22680 21728 0 net25
rlabel metal3 118706 111496 118706 111496 0 net250
rlabel metal3 1302 84168 1302 84168 0 net251
rlabel metal3 1302 48552 1302 48552 0 net252
rlabel metal2 37128 2030 37128 2030 0 net253
rlabel metal2 118104 96600 118104 96600 0 net254
rlabel metal2 118104 46648 118104 46648 0 net255
rlabel metal2 118104 2744 118104 2744 0 net256
rlabel metal3 118720 16968 118720 16968 0 net257
rlabel metal3 1302 6888 1302 6888 0 net258
rlabel metal3 1302 107688 1302 107688 0 net259
rlabel metal3 35896 101752 35896 101752 0 net26
rlabel metal3 1302 54600 1302 54600 0 net260
rlabel metal2 118104 101304 118104 101304 0 net261
rlabel metal2 49896 2590 49896 2590 0 net262
rlabel metal2 19040 116312 19040 116312 0 net263
rlabel metal2 109704 2030 109704 2030 0 net264
rlabel metal3 1302 85512 1302 85512 0 net265
rlabel metal2 27720 2030 27720 2030 0 net266
rlabel metal2 109032 2030 109032 2030 0 net267
rlabel metal3 69216 115864 69216 115864 0 net268
rlabel metal2 41888 115864 41888 115864 0 net269
rlabel metal3 45920 105784 45920 105784 0 net27
rlabel metal3 2758 115752 2758 115752 0 net270
rlabel metal2 86912 114744 86912 114744 0 net271
rlabel metal2 94304 116312 94304 116312 0 net272
rlabel metal2 51352 116704 51352 116704 0 net273
rlabel metal3 1302 16968 1302 16968 0 net274
rlabel metal3 118706 70728 118706 70728 0 net275
rlabel metal2 118104 82600 118104 82600 0 net276
rlabel metal3 118706 106792 118706 106792 0 net277
rlabel metal3 1302 109704 1302 109704 0 net278
rlabel metal2 97944 117040 97944 117040 0 net279
rlabel metal3 71624 26040 71624 26040 0 net28
rlabel metal2 32424 798 32424 798 0 net280
rlabel metal2 104328 1246 104328 1246 0 net281
rlabel metal3 1302 18312 1302 18312 0 net282
rlabel metal2 43176 117810 43176 117810 0 net283
rlabel metal2 75432 2030 75432 2030 0 net284
rlabel metal3 118706 56616 118706 56616 0 net285
rlabel metal2 26936 3640 26936 3640 0 net29
rlabel metal3 39928 115528 39928 115528 0 net3
rlabel metal2 101864 49336 101864 49336 0 net30
rlabel metal2 68040 67200 68040 67200 0 net31
rlabel metal3 106232 115528 106232 115528 0 net32
rlabel metal2 3360 4200 3360 4200 0 net33
rlabel metal2 3360 116536 3360 116536 0 net34
rlabel metal2 63784 3696 63784 3696 0 net35
rlabel metal2 3304 52136 3304 52136 0 net36
rlabel metal2 32200 63000 32200 63000 0 net37
rlabel metal2 3360 35000 3360 35000 0 net38
rlabel metal2 44520 88844 44520 88844 0 net39
rlabel metal2 51240 116480 51240 116480 0 net4
rlabel metal2 26040 67760 26040 67760 0 net40
rlabel metal3 54376 44968 54376 44968 0 net41
rlabel metal2 3304 60144 3304 60144 0 net42
rlabel metal2 96376 4760 96376 4760 0 net43
rlabel metal2 46088 5152 46088 5152 0 net44
rlabel metal2 24360 74816 24360 74816 0 net45
rlabel metal2 108360 58912 108360 58912 0 net46
rlabel metal2 83272 70392 83272 70392 0 net47
rlabel metal2 93016 29456 93016 29456 0 net48
rlabel metal2 43624 116144 43624 116144 0 net49
rlabel metal3 73080 63280 73080 63280 0 net5
rlabel metal2 114968 5880 114968 5880 0 net50
rlabel metal3 80696 116536 80696 116536 0 net51
rlabel metal2 114856 61880 114856 61880 0 net52
rlabel metal2 91952 20160 91952 20160 0 net53
rlabel metal2 91560 58016 91560 58016 0 net54
rlabel metal2 101864 26208 101864 26208 0 net55
rlabel metal3 70224 56840 70224 56840 0 net56
rlabel metal3 109984 3640 109984 3640 0 net57
rlabel metal2 33544 57512 33544 57512 0 net58
rlabel metal2 24360 29344 24360 29344 0 net59
rlabel metal2 43232 4648 43232 4648 0 net6
rlabel metal2 76664 57288 76664 57288 0 net60
rlabel metal2 62216 72968 62216 72968 0 net61
rlabel metal2 31080 27888 31080 27888 0 net62
rlabel metal2 115528 4704 115528 4704 0 net63
rlabel metal2 26040 39760 26040 39760 0 net64
rlabel metal2 24024 116536 24024 116536 0 net65
rlabel metal3 39032 99400 39032 99400 0 net66
rlabel metal2 100072 78288 100072 78288 0 net67
rlabel metal3 30632 93016 30632 93016 0 net68
rlabel metal2 22680 82376 22680 82376 0 net69
rlabel metal3 60032 3640 60032 3640 0 net7
rlabel metal3 9632 97720 9632 97720 0 net70
rlabel metal3 6692 3640 6692 3640 0 net71
rlabel metal2 3304 25648 3304 25648 0 net72
rlabel metal4 73304 63224 73304 63224 0 net73
rlabel metal3 70224 25816 70224 25816 0 net74
rlabel metal2 78680 61320 78680 61320 0 net75
rlabel metal2 101640 85400 101640 85400 0 net76
rlabel metal2 7560 93128 7560 93128 0 net77
rlabel metal2 29400 28784 29400 28784 0 net78
rlabel metal2 3304 30240 3304 30240 0 net79
rlabel metal2 22680 49000 22680 49000 0 net8
rlabel metal3 116984 116536 116984 116536 0 net80
rlabel metal2 3360 71624 3360 71624 0 net81
rlabel metal3 101528 94584 101528 94584 0 net82
rlabel metal2 115192 42560 115192 42560 0 net83
rlabel metal3 77784 27720 77784 27720 0 net84
rlabel metal2 99848 110880 99848 110880 0 net85
rlabel metal2 30408 84504 30408 84504 0 net86
rlabel metal3 42448 48776 42448 48776 0 net87
rlabel metal3 109928 74200 109928 74200 0 net88
rlabel metal2 98392 4256 98392 4256 0 net89
rlabel metal3 111552 35224 111552 35224 0 net9
rlabel metal2 114856 37184 114856 37184 0 net90
rlabel metal2 3360 63784 3360 63784 0 net91
rlabel metal2 114800 5208 114800 5208 0 net92
rlabel metal2 20664 3696 20664 3696 0 net93
rlabel metal2 60088 42112 60088 42112 0 net94
rlabel metal2 108248 49672 108248 49672 0 net95
rlabel metal2 95928 116480 95928 116480 0 net96
rlabel metal3 78960 60256 78960 60256 0 net97
rlabel metal2 98280 34272 98280 34272 0 net98
rlabel metal2 29400 81704 29400 81704 0 net99
rlabel metal3 117250 21000 117250 21000 0 wb_clk_i
rlabel metal2 22064 116536 22064 116536 0 wb_rst_i
rlabel metal3 117586 41832 117586 41832 0 wbs_ack_o
rlabel metal2 38192 116536 38192 116536 0 wbs_cyc_i
rlabel metal2 116872 104440 116872 104440 0 wbs_dat_i[0]
rlabel metal3 1358 92792 1358 92792 0 wbs_dat_i[10]
rlabel metal3 1582 101640 1582 101640 0 wbs_dat_i[11]
rlabel metal3 1246 96936 1246 96936 0 wbs_dat_i[12]
rlabel metal2 3864 4592 3864 4592 0 wbs_dat_i[13]
rlabel metal2 1960 25200 1960 25200 0 wbs_dat_i[14]
rlabel metal2 117096 62776 117096 62776 0 wbs_dat_i[15]
rlabel metal2 69104 3416 69104 3416 0 wbs_dat_i[16]
rlabel metal2 81872 115864 81872 115864 0 wbs_dat_i[17]
rlabel metal2 110936 117936 110936 117936 0 wbs_dat_i[18]
rlabel metal2 5936 116536 5936 116536 0 wbs_dat_i[19]
rlabel metal2 18032 4200 18032 4200 0 wbs_dat_i[1]
rlabel metal3 1302 29624 1302 29624 0 wbs_dat_i[20]
rlabel metal2 114856 117922 114856 117922 0 wbs_dat_i[21]
rlabel metal2 1848 71120 1848 71120 0 wbs_dat_i[22]
rlabel metal3 118202 94248 118202 94248 0 wbs_dat_i[23]
rlabel metal3 118202 39704 118202 39704 0 wbs_dat_i[24]
rlabel metal2 83496 2086 83496 2086 0 wbs_dat_i[25]
rlabel metal2 99288 116536 99288 116536 0 wbs_dat_i[26]
rlabel metal2 28784 115864 28784 115864 0 wbs_dat_i[27]
rlabel metal2 37912 3416 37912 3416 0 wbs_dat_i[28]
rlabel metal2 117096 73696 117096 73696 0 wbs_dat_i[29]
rlabel metal2 98000 4200 98000 4200 0 wbs_dat_i[2]
rlabel metal2 117096 36008 117096 36008 0 wbs_dat_i[30]
rlabel metal2 1960 63672 1960 63672 0 wbs_dat_i[31]
rlabel metal3 118202 4872 118202 4872 0 wbs_dat_i[3]
rlabel metal2 21560 4032 21560 4032 0 wbs_dat_i[4]
rlabel metal2 59864 2926 59864 2926 0 wbs_dat_i[5]
rlabel metal2 116872 52696 116872 52696 0 wbs_dat_i[6]
rlabel metal2 95144 116928 95144 116928 0 wbs_dat_i[7]
rlabel metal3 118090 107688 118090 107688 0 wbs_dat_i[8]
rlabel metal2 116200 6384 116200 6384 0 wbs_dat_i[9]
rlabel metal3 1358 24360 1358 24360 0 wbs_dat_o[0]
rlabel metal3 117586 68712 117586 68712 0 wbs_dat_o[10]
rlabel metal2 2184 2478 2184 2478 0 wbs_dat_o[11]
rlabel metal3 117586 110376 117586 110376 0 wbs_dat_o[12]
rlabel metal3 91784 116536 91784 116536 0 wbs_dat_o[13]
rlabel metal3 117586 14280 117586 14280 0 wbs_dat_o[14]
rlabel metal2 86968 115696 86968 115696 0 wbs_dat_o[15]
rlabel metal3 1358 33768 1358 33768 0 wbs_dat_o[16]
rlabel metal3 1358 37800 1358 37800 0 wbs_dat_o[17]
rlabel metal2 80808 798 80808 798 0 wbs_dat_o[18]
rlabel metal2 168 2198 168 2198 0 wbs_dat_o[19]
rlabel metal2 94920 798 94920 798 0 wbs_dat_o[1]
rlabel metal3 1358 56616 1358 56616 0 wbs_dat_o[20]
rlabel metal3 1358 104328 1358 104328 0 wbs_dat_o[21]
rlabel metal2 32088 116480 32088 116480 0 wbs_dat_o[22]
rlabel metal3 1358 39144 1358 39144 0 wbs_dat_o[23]
rlabel metal2 25032 2926 25032 2926 0 wbs_dat_o[24]
rlabel metal2 8904 2086 8904 2086 0 wbs_dat_o[25]
rlabel metal2 62664 117530 62664 117530 0 wbs_dat_o[26]
rlabel metal2 35112 117530 35112 117530 0 wbs_dat_o[27]
rlabel metal2 64680 798 64680 798 0 wbs_dat_o[28]
rlabel metal3 84168 116536 84168 116536 0 wbs_dat_o[29]
rlabel metal2 115528 33544 115528 33544 0 wbs_dat_o[2]
rlabel metal3 1358 78680 1358 78680 0 wbs_dat_o[30]
rlabel metal3 117586 92904 117586 92904 0 wbs_dat_o[31]
rlabel metal2 26376 2478 26376 2478 0 wbs_dat_o[3]
rlabel metal2 46536 798 46536 798 0 wbs_dat_o[4]
rlabel metal3 1358 10248 1358 10248 0 wbs_dat_o[5]
rlabel metal2 115416 89712 115416 89712 0 wbs_dat_o[6]
rlabel metal2 72744 2478 72744 2478 0 wbs_dat_o[7]
rlabel metal2 78792 117530 78792 117530 0 wbs_dat_o[8]
rlabel metal2 78120 117922 78120 117922 0 wbs_dat_o[9]
rlabel metal3 1246 111048 1246 111048 0 wbs_sel_i[0]
rlabel metal2 12824 117922 12824 117922 0 wbs_sel_i[1]
rlabel metal2 86576 4200 86576 4200 0 wbs_sel_i[2]
rlabel metal3 1246 26376 1246 26376 0 wbs_sel_i[3]
rlabel metal2 1848 99344 1848 99344 0 wbs_stb_i
rlabel metal2 115864 59528 115864 59528 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 120000 120000
<< end >>
